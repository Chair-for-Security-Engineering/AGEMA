module Reg1(x, y);
 input [133:0] x;
 output [132:0] y;

  assign y[0] = x[133];
  assign y[5] = x[0];
  assign y[6] = x[11];
  assign y[7] = x[22];
  assign y[8] = x[33];
  assign y[9] = x[44];
  assign y[10] = x[55];
  assign y[11] = x[60];
  assign y[12] = x[61];
  assign y[13] = x[62];
  assign y[14] = x[63];
  assign y[15] = x[1];
  assign y[16] = x[2];
  assign y[17] = x[3];
  assign y[18] = x[4];
  assign y[19] = x[5];
  assign y[20] = x[6];
  assign y[21] = x[7];
  assign y[22] = x[8];
  assign y[23] = x[9];
  assign y[24] = x[10];
  assign y[25] = x[12];
  assign y[26] = x[13];
  assign y[27] = x[14];
  assign y[28] = x[15];
  assign y[29] = x[16];
  assign y[30] = x[17];
  assign y[31] = x[18];
  assign y[32] = x[19];
  assign y[33] = x[20];
  assign y[34] = x[21];
  assign y[35] = x[23];
  assign y[36] = x[24];
  assign y[37] = x[25];
  assign y[38] = x[26];
  assign y[39] = x[27];
  assign y[40] = x[28];
  assign y[41] = x[29];
  assign y[42] = x[30];
  assign y[43] = x[31];
  assign y[44] = x[32];
  assign y[45] = x[34];
  assign y[46] = x[35];
  assign y[47] = x[36];
  assign y[48] = x[37];
  assign y[49] = x[38];
  assign y[50] = x[39];
  assign y[51] = x[40];
  assign y[52] = x[41];
  assign y[53] = x[42];
  assign y[54] = x[43];
  assign y[55] = x[45];
  assign y[56] = x[46];
  assign y[57] = x[47];
  assign y[58] = x[48];
  assign y[59] = x[49];
  assign y[60] = x[50];
  assign y[61] = x[51];
  assign y[62] = x[52];
  assign y[63] = x[53];
  assign y[64] = x[54];
  assign y[65] = x[56];
  assign y[66] = x[57];
  assign y[67] = x[58];
  assign y[68] = x[59];
  register_stage #(.WIDTH(68)) inst_0(.clk(x[128]), .D({x[129],x[130],x[131],x[132],x[64],x[75],x[86],x[97],x[108],x[119],x[124],x[125],x[126],x[127],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[120],x[121],x[122],x[123]}), .Q({y[1],y[2],y[3],y[4],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132]}));
endmodule

module Reg2(x, y);
 input [185:0] x;
 output [184:0] y;

  assign y[0] = x[181];
  assign y[1] = x[182];
  assign y[2] = x[183];
  assign y[3] = x[184];
  assign y[4] = x[185];
  assign y[25] = x[0];
  assign y[26] = x[1];
  assign y[27] = x[2];
  assign y[28] = x[3];
  assign y[29] = x[4];
  assign y[30] = x[55];
  assign y[31] = x[56];
  assign y[32] = x[57];
  assign y[33] = x[58];
  assign y[34] = x[59];
  assign y[35] = x[75];
  assign y[36] = x[76];
  assign y[37] = x[77];
  assign y[38] = x[78];
  assign y[39] = x[79];
  assign y[40] = x[5];
  assign y[41] = x[6];
  assign y[42] = x[7];
  assign y[43] = x[8];
  assign y[44] = x[9];
  assign y[45] = x[10];
  assign y[46] = x[11];
  assign y[47] = x[12];
  assign y[48] = x[13];
  assign y[49] = x[14];
  assign y[50] = x[15];
  assign y[51] = x[16];
  assign y[52] = x[17];
  assign y[53] = x[18];
  assign y[54] = x[19];
  assign y[55] = x[20];
  assign y[56] = x[21];
  assign y[57] = x[22];
  assign y[58] = x[23];
  assign y[59] = x[24];
  assign y[60] = x[25];
  assign y[61] = x[26];
  assign y[62] = x[27];
  assign y[63] = x[28];
  assign y[64] = x[29];
  assign y[65] = x[30];
  assign y[66] = x[31];
  assign y[67] = x[32];
  assign y[68] = x[33];
  assign y[69] = x[34];
  assign y[70] = x[35];
  assign y[71] = x[36];
  assign y[72] = x[37];
  assign y[73] = x[38];
  assign y[74] = x[39];
  assign y[75] = x[40];
  assign y[76] = x[41];
  assign y[77] = x[42];
  assign y[78] = x[43];
  assign y[79] = x[44];
  assign y[80] = x[45];
  assign y[81] = x[46];
  assign y[82] = x[47];
  assign y[83] = x[48];
  assign y[84] = x[49];
  assign y[85] = x[50];
  assign y[86] = x[51];
  assign y[87] = x[52];
  assign y[88] = x[53];
  assign y[89] = x[54];
  assign y[90] = x[60];
  assign y[91] = x[61];
  assign y[92] = x[62];
  assign y[93] = x[63];
  assign y[94] = x[64];
  assign y[95] = x[65];
  assign y[96] = x[66];
  assign y[97] = x[67];
  assign y[98] = x[68];
  assign y[99] = x[69];
  assign y[100] = x[70];
  assign y[101] = x[71];
  assign y[102] = x[72];
  assign y[103] = x[73];
  assign y[104] = x[74];
  register_stage #(.WIDTH(100)) inst_0(.clk(x[160]), .D({x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[80],x[81],x[82],x[83],x[84],x[135],x[136],x[137],x[138],x[139],x[155],x[156],x[157],x[158],x[159],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154]}), .Q({y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [302:0] x;
 output [169:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx4 Fx4_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx5 Fx5_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx9 Fx9_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx10 Fx10_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx14 Fx14_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx15 Fx15_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx19 Fx19_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx20 Fx20_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx24 Fx24_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx25 Fx25_inst(.x({x[19], x[18], x[17], x[16], x[15]}), .y(y[10]));
  Fx26 Fx26_inst(.x({x[20], x[18]}), .y(y[11]));
  Fx27 Fx27_inst(.x({x[21], x[17]}), .y(y[12]));
  Fx28 Fx28_inst(.x({x[22], x[16]}), .y(y[13]));
  Fx29 Fx29_inst(.x({x[23], x[15]}), .y(y[14]));
  Fx30 Fx30_inst(.x({x[28], x[27], x[26], x[25], x[24]}), .y(y[15]));
  Fx31 Fx31_inst(.x({x[29], x[27]}), .y(y[16]));
  Fx32 Fx32_inst(.x({x[30], x[26]}), .y(y[17]));
  Fx33 Fx33_inst(.x({x[31], x[25]}), .y(y[18]));
  Fx34 Fx34_inst(.x({x[32], x[24]}), .y(y[19]));
  Fx35 Fx35_inst(.x({x[37], x[36], x[35], x[34], x[33]}), .y(y[20]));
  Fx36 Fx36_inst(.x({x[38], x[36]}), .y(y[21]));
  Fx37 Fx37_inst(.x({x[39], x[35]}), .y(y[22]));
  Fx38 Fx38_inst(.x({x[40], x[34]}), .y(y[23]));
  Fx39 Fx39_inst(.x({x[41], x[33]}), .y(y[24]));
  Fx40 Fx40_inst(.x({x[46], x[45], x[44], x[43], x[42]}), .y(y[25]));
  Fx41 Fx41_inst(.x({x[47], x[45]}), .y(y[26]));
  Fx42 Fx42_inst(.x({x[48], x[44]}), .y(y[27]));
  Fx43 Fx43_inst(.x({x[49], x[43]}), .y(y[28]));
  Fx44 Fx44_inst(.x({x[50], x[42]}), .y(y[29]));
  Fx45 Fx45_inst(.x({x[55], x[54], x[53], x[52], x[51]}), .y(y[30]));
  Fx46 Fx46_inst(.x({x[56], x[54]}), .y(y[31]));
  Fx47 Fx47_inst(.x({x[57], x[53]}), .y(y[32]));
  Fx48 Fx48_inst(.x({x[58], x[52]}), .y(y[33]));
  Fx49 Fx49_inst(.x({x[59], x[51]}), .y(y[34]));
  Fx50 Fx50_inst(.x({x[64], x[63], x[62], x[61], x[60]}), .y(y[35]));
  Fx51 Fx51_inst(.x({x[65], x[63]}), .y(y[36]));
  Fx52 Fx52_inst(.x({x[66], x[62]}), .y(y[37]));
  Fx53 Fx53_inst(.x({x[67], x[61]}), .y(y[38]));
  Fx54 Fx54_inst(.x({x[68], x[60]}), .y(y[39]));
  Fx55 Fx55_inst(.x({x[73], x[72], x[71], x[70], x[69]}), .y(y[40]));
  Fx56 Fx56_inst(.x({x[74], x[72]}), .y(y[41]));
  Fx57 Fx57_inst(.x({x[75], x[71]}), .y(y[42]));
  Fx58 Fx58_inst(.x({x[76], x[70]}), .y(y[43]));
  Fx59 Fx59_inst(.x({x[77], x[69]}), .y(y[44]));
  Fx60 Fx60_inst(.x({x[82], x[81], x[80], x[79], x[78]}), .y(y[45]));
  Fx61 Fx61_inst(.x({x[83], x[81]}), .y(y[46]));
  Fx62 Fx62_inst(.x({x[84], x[80]}), .y(y[47]));
  Fx63 Fx63_inst(.x({x[85], x[79]}), .y(y[48]));
  Fx64 Fx64_inst(.x({x[86], x[78]}), .y(y[49]));
  Fx65 Fx65_inst(.x({x[91], x[90], x[89], x[88], x[87]}), .y(y[50]));
  Fx66 Fx66_inst(.x({x[92], x[90]}), .y(y[51]));
  Fx67 Fx67_inst(.x({x[93], x[89]}), .y(y[52]));
  Fx68 Fx68_inst(.x({x[94], x[88]}), .y(y[53]));
  Fx69 Fx69_inst(.x({x[95], x[87]}), .y(y[54]));
  Fx70 Fx70_inst(.x({x[100], x[99], x[98], x[97], x[96]}), .y(y[55]));
  Fx71 Fx71_inst(.x({x[101], x[99]}), .y(y[56]));
  Fx72 Fx72_inst(.x({x[102], x[98]}), .y(y[57]));
  Fx73 Fx73_inst(.x({x[103], x[97]}), .y(y[58]));
  Fx74 Fx74_inst(.x({x[104], x[96]}), .y(y[59]));
  Fx75 Fx75_inst(.x({x[109], x[108], x[107], x[106], x[105]}), .y(y[60]));
  Fx76 Fx76_inst(.x({x[110], x[108]}), .y(y[61]));
  Fx77 Fx77_inst(.x({x[111], x[107]}), .y(y[62]));
  Fx78 Fx78_inst(.x({x[112], x[106]}), .y(y[63]));
  Fx79 Fx79_inst(.x({x[113], x[105]}), .y(y[64]));
  Fx80 Fx80_inst(.x({x[118], x[117], x[116], x[115], x[114]}), .y(y[65]));
  Fx81 Fx81_inst(.x({x[119], x[117]}), .y(y[66]));
  Fx82 Fx82_inst(.x({x[120], x[116]}), .y(y[67]));
  Fx83 Fx83_inst(.x({x[121], x[115]}), .y(y[68]));
  Fx84 Fx84_inst(.x({x[122], x[114]}), .y(y[69]));
  Fx85 Fx85_inst(.x({x[127], x[126], x[125], x[124], x[123]}), .y(y[70]));
  Fx86 Fx86_inst(.x({x[128], x[126]}), .y(y[71]));
  Fx87 Fx87_inst(.x({x[129], x[125]}), .y(y[72]));
  Fx88 Fx88_inst(.x({x[130], x[124]}), .y(y[73]));
  Fx89 Fx89_inst(.x({x[131], x[123]}), .y(y[74]));
  Fx90 Fx90_inst(.x({x[136], x[135], x[134], x[133], x[132]}), .y(y[75]));
  Fx91 Fx91_inst(.x({x[137], x[135]}), .y(y[76]));
  Fx92 Fx92_inst(.x({x[138], x[134]}), .y(y[77]));
  Fx93 Fx93_inst(.x({x[139], x[133]}), .y(y[78]));
  Fx94 Fx94_inst(.x({x[140], x[132]}), .y(y[79]));
  Fx95 Fx95_inst(.x({x[145], x[144], x[143], x[142], x[141]}), .y(y[80]));
  Fx96 Fx96_inst(.x({x[146], x[144]}), .y(y[81]));
  Fx97 Fx97_inst(.x({x[147], x[143]}), .y(y[82]));
  Fx98 Fx98_inst(.x({x[148], x[142]}), .y(y[83]));
  Fx99 Fx99_inst(.x({x[149], x[141]}), .y(y[84]));
  Fx100 Fx100_inst(.x({x[154], x[153], x[152], x[151], x[150]}), .y(y[85]));
  Fx101 Fx101_inst(.x({x[155], x[153]}), .y(y[86]));
  Fx102 Fx102_inst(.x({x[156], x[152]}), .y(y[87]));
  Fx103 Fx103_inst(.x({x[157], x[151]}), .y(y[88]));
  Fx104 Fx104_inst(.x({x[158], x[150]}), .y(y[89]));
  Fx105 Fx105_inst(.x({x[163], x[162], x[161], x[160], x[159]}), .y(y[90]));
  Fx106 Fx106_inst(.x({x[164], x[162]}), .y(y[91]));
  Fx107 Fx107_inst(.x({x[165], x[161]}), .y(y[92]));
  Fx108 Fx108_inst(.x({x[166], x[160]}), .y(y[93]));
  Fx109 Fx109_inst(.x({x[167], x[159]}), .y(y[94]));
  Fx110 Fx110_inst(.x({x[172], x[171], x[170], x[169], x[168]}), .y(y[95]));
  Fx111 Fx111_inst(.x({x[173], x[171]}), .y(y[96]));
  Fx112 Fx112_inst(.x({x[174], x[170]}), .y(y[97]));
  Fx113 Fx113_inst(.x({x[175], x[169]}), .y(y[98]));
  Fx114 Fx114_inst(.x({x[176], x[168]}), .y(y[99]));
  Fx115 Fx115_inst(.x({x[181], x[180], x[179], x[178], x[177]}), .y(y[100]));
  Fx116 Fx116_inst(.x({x[182], x[180]}), .y(y[101]));
  Fx117 Fx117_inst(.x({x[183], x[179]}), .y(y[102]));
  Fx118 Fx118_inst(.x({x[184], x[178]}), .y(y[103]));
  Fx119 Fx119_inst(.x({x[185], x[177]}), .y(y[104]));
  Fx120 Fx120_inst(.x({x[190], x[189], x[188], x[187], x[186]}), .y(y[105]));
  Fx121 Fx121_inst(.x({x[191], x[189]}), .y(y[106]));
  Fx122 Fx122_inst(.x({x[192], x[188]}), .y(y[107]));
  Fx123 Fx123_inst(.x({x[193], x[187]}), .y(y[108]));
  Fx124 Fx124_inst(.x({x[194], x[186]}), .y(y[109]));
  Fx125 Fx125_inst(.x({x[199], x[198], x[197], x[196], x[195]}), .y(y[110]));
  Fx126 Fx126_inst(.x({x[200], x[198]}), .y(y[111]));
  Fx127 Fx127_inst(.x({x[201], x[197]}), .y(y[112]));
  Fx128 Fx128_inst(.x({x[202], x[196]}), .y(y[113]));
  Fx129 Fx129_inst(.x({x[203], x[195]}), .y(y[114]));
  Fx130 Fx130_inst(.x({x[208], x[207], x[206], x[205], x[204]}), .y(y[115]));
  Fx131 Fx131_inst(.x({x[209], x[207]}), .y(y[116]));
  Fx132 Fx132_inst(.x({x[210], x[206]}), .y(y[117]));
  Fx133 Fx133_inst(.x({x[211], x[205]}), .y(y[118]));
  Fx134 Fx134_inst(.x({x[212], x[204]}), .y(y[119]));
  Fx135 Fx135_inst(.x({x[217], x[216], x[215], x[214], x[213]}), .y(y[120]));
  Fx136 Fx136_inst(.x({x[218], x[216]}), .y(y[121]));
  Fx137 Fx137_inst(.x({x[219], x[215]}), .y(y[122]));
  Fx138 Fx138_inst(.x({x[220], x[214]}), .y(y[123]));
  Fx139 Fx139_inst(.x({x[221], x[213]}), .y(y[124]));
  Fx140 Fx140_inst(.x({x[226], x[225], x[224], x[223], x[222]}), .y(y[125]));
  Fx141 Fx141_inst(.x({x[227], x[225]}), .y(y[126]));
  Fx142 Fx142_inst(.x({x[228], x[224]}), .y(y[127]));
  Fx143 Fx143_inst(.x({x[229], x[223]}), .y(y[128]));
  Fx144 Fx144_inst(.x({x[230], x[222]}), .y(y[129]));
  Fx145 Fx145_inst(.x({x[235], x[234], x[233], x[232], x[231]}), .y(y[130]));
  Fx146 Fx146_inst(.x({x[236], x[234]}), .y(y[131]));
  Fx147 Fx147_inst(.x({x[237], x[233]}), .y(y[132]));
  Fx148 Fx148_inst(.x({x[238], x[232]}), .y(y[133]));
  Fx149 Fx149_inst(.x({x[239], x[231]}), .y(y[134]));
  Fx150 Fx150_inst(.x({x[244], x[243], x[242], x[241], x[240]}), .y(y[135]));
  Fx151 Fx151_inst(.x({x[245], x[243]}), .y(y[136]));
  Fx152 Fx152_inst(.x({x[246], x[242]}), .y(y[137]));
  Fx153 Fx153_inst(.x({x[247], x[241]}), .y(y[138]));
  Fx154 Fx154_inst(.x({x[248], x[240]}), .y(y[139]));
  Fx155 Fx155_inst(.x({x[253], x[252], x[251], x[250], x[249]}), .y(y[140]));
  Fx156 Fx156_inst(.x({x[254], x[252]}), .y(y[141]));
  Fx157 Fx157_inst(.x({x[255], x[251]}), .y(y[142]));
  Fx158 Fx158_inst(.x({x[256], x[250]}), .y(y[143]));
  Fx159 Fx159_inst(.x({x[257], x[249]}), .y(y[144]));
  Fx160 Fx160_inst(.x({x[262], x[261], x[260], x[259], x[258]}), .y(y[145]));
  Fx161 Fx161_inst(.x({x[263], x[261]}), .y(y[146]));
  Fx162 Fx162_inst(.x({x[264], x[260]}), .y(y[147]));
  Fx163 Fx163_inst(.x({x[265], x[259]}), .y(y[148]));
  Fx164 Fx164_inst(.x({x[266], x[258]}), .y(y[149]));
  Fx165 Fx165_inst(.x({x[271], x[270], x[269], x[268], x[267]}), .y(y[150]));
  Fx166 Fx166_inst(.x({x[272], x[270]}), .y(y[151]));
  Fx167 Fx167_inst(.x({x[273], x[269]}), .y(y[152]));
  Fx168 Fx168_inst(.x({x[274], x[268]}), .y(y[153]));
  Fx169 Fx169_inst(.x({x[275], x[267]}), .y(y[154]));
  Fx170 Fx170_inst(.x({x[280], x[279], x[278], x[277], x[276]}), .y(y[155]));
  Fx171 Fx171_inst(.x({x[281], x[279]}), .y(y[156]));
  Fx172 Fx172_inst(.x({x[282], x[278]}), .y(y[157]));
  Fx173 Fx173_inst(.x({x[283], x[277]}), .y(y[158]));
  Fx174 Fx174_inst(.x({x[284], x[276]}), .y(y[159]));
  Fx175 Fx175_inst(.x({x[289], x[288], x[287], x[286], x[285]}), .y(y[160]));
  Fx176 Fx176_inst(.x({x[290], x[288]}), .y(y[161]));
  Fx177 Fx177_inst(.x({x[291], x[287]}), .y(y[162]));
  Fx178 Fx178_inst(.x({x[292], x[286]}), .y(y[163]));
  Fx179 Fx179_inst(.x({x[293], x[285]}), .y(y[164]));
  Fx180 Fx180_inst(.x({x[298], x[297], x[296], x[295], x[294]}), .y(y[165]));
  Fx181 Fx181_inst(.x({x[299], x[297]}), .y(y[166]));
  Fx182 Fx182_inst(.x({x[300], x[296]}), .y(y[167]));
  Fx183 Fx183_inst(.x({x[301], x[295]}), .y(y[168]));
  Fx184 Fx184_inst(.x({x[302], x[294]}), .y(y[169]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind66(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind67(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind68(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind69(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind70(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind71(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind72(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind73(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind74(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind75(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind76(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind77(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind78(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind79(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind80(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind81(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind82(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind83(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind84(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind85(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind86(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind87(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind88(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind89(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind90(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind91(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind92(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind93(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind94(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind95(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind96(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind97(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind98(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind99(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind100(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind101(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind102(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind103(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind104(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind105(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind106(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind107(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind108(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind109(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind110(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind111(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind112(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind113(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind114(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind115(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind116(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind117(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind118(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind119(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind120(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind121(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind122(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind123(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind124(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind125(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[8];
  assign t[11] = t[15] ^ x[10];
  assign t[12] = (x[2] & x[3]);
  assign t[13] = (x[2] & x[5]);
  assign t[14] = (x[2] & x[7]);
  assign t[15] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = t[6] | t[8];
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[7] | t[4]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = t[0] ^ t[1];
endmodule

module R1ind126(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6] & t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[11] & t[10]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind127(x, y);
 input [8:0] x;
 output y;

 wire [12:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = (x[2] & x[3]);
  assign t[11] = (x[2] & x[5]);
  assign t[12] = (x[2] & x[7]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[9] & t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = t[10] ^ x[4];
  assign t[8] = t[11] ^ x[6];
  assign t[9] = t[12] ^ x[8];
  assign y = t[0] ^ t[1];
endmodule

module R1ind128(x, y);
 input [10:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = x[0] ^ x[1];
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[10];
  assign t[13] = (x[2] & x[3]);
  assign t[14] = (x[2] & x[5]);
  assign t[15] = (x[2] & x[7]);
  assign t[16] = (x[2] & x[9]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[9] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[12]);
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = t[13] ^ x[4];
  assign y = t[0] ^ t[1];
endmodule

module R1ind129(x, y);
 input [11:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[2] = t[6] ^ x[2];
  assign t[3] = t[7] ^ x[5];
  assign t[4] = t[8] ^ x[8];
  assign t[5] = t[9] ^ x[11];
  assign t[6] = (x[0] & x[1]);
  assign t[7] = (x[3] & x[4]);
  assign t[8] = (x[6] & x[7]);
  assign t[9] = (x[9] & x[10]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind130(x, y);
 input [79:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = (x[11] & x[12]);
  assign t[101] = (x[14] & x[15]);
  assign t[102] = (x[17] & x[18]);
  assign t[103] = (x[20] & x[21]);
  assign t[104] = (x[20] & x[25]);
  assign t[105] = (x[20] & x[27]);
  assign t[106] = (x[29] & x[30]);
  assign t[107] = (x[32] & x[33]);
  assign t[108] = (x[37] & x[38]);
  assign t[109] = (x[20] & x[42]);
  assign t[10] = ~(x[3]);
  assign t[110] = (x[29] & x[44]);
  assign t[111] = (x[29] & x[46]);
  assign t[112] = (x[32] & x[48]);
  assign t[113] = (x[32] & x[50]);
  assign t[114] = (x[52] & x[53]);
  assign t[115] = (x[37] & x[55]);
  assign t[116] = (x[37] & x[57]);
  assign t[117] = (x[59] & x[60]);
  assign t[118] = (x[29] & x[62]);
  assign t[119] = (x[32] & x[64]);
  assign t[11] = t[16] ? x[7] : x[6];
  assign t[120] = (x[52] & x[66]);
  assign t[121] = (x[52] & x[68]);
  assign t[122] = (x[37] & x[70]);
  assign t[123] = (x[59] & x[72]);
  assign t[124] = (x[59] & x[74]);
  assign t[125] = (x[52] & x[76]);
  assign t[126] = (x[59] & x[78]);
  assign t[12] = x[4] ? t[18] : t[17];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[14] = ~(t[70] & t[71]);
  assign t[15] = ~(t[72] & t[73]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = t[24] ^ t[25];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = x[4] ? t[29] : t[28];
  assign t[21] = ~(t[72]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = t[32] | t[74];
  assign t[24] = t[16] ? x[24] : x[23];
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = ~(t[35] & t[36]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[75]);
  assign t[31] = ~(t[76]);
  assign t[32] = ~(t[43] | t[30]);
  assign t[33] = ~(t[44] & t[45]);
  assign t[34] = t[46] | t[77];
  assign t[35] = ~(t[47] & t[48]);
  assign t[36] = t[49] | t[78];
  assign t[37] = t[50] ? x[36] : x[35];
  assign t[38] = ~(t[51] & t[52]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[55] | t[79];
  assign t[41] = t[16] ? x[41] : x[40];
  assign t[42] = ~(t[56] & t[57]);
  assign t[43] = ~(t[80]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[82]);
  assign t[46] = ~(t[58] | t[44]);
  assign t[47] = ~(t[83]);
  assign t[48] = ~(t[84]);
  assign t[49] = ~(t[59] | t[47]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[21]);
  assign t[51] = ~(t[60] & t[61]);
  assign t[52] = t[62] | t[85];
  assign t[53] = ~(t[86]);
  assign t[54] = ~(t[87]);
  assign t[55] = ~(t[63] | t[53]);
  assign t[56] = ~(t[64] & t[65]);
  assign t[57] = t[66] | t[88];
  assign t[58] = ~(t[89]);
  assign t[59] = ~(t[90]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[91]);
  assign t[61] = ~(t[92]);
  assign t[62] = ~(t[67] | t[60]);
  assign t[63] = ~(t[93]);
  assign t[64] = ~(t[94]);
  assign t[65] = ~(t[95]);
  assign t[66] = ~(t[68] | t[64]);
  assign t[67] = ~(t[96]);
  assign t[68] = ~(t[97]);
  assign t[69] = t[98] ^ x[2];
  assign t[6] = t[11] ^ t[7];
  assign t[70] = t[99] ^ x[10];
  assign t[71] = t[100] ^ x[13];
  assign t[72] = t[101] ^ x[16];
  assign t[73] = t[102] ^ x[19];
  assign t[74] = t[103] ^ x[22];
  assign t[75] = t[104] ^ x[26];
  assign t[76] = t[105] ^ x[28];
  assign t[77] = t[106] ^ x[31];
  assign t[78] = t[107] ^ x[34];
  assign t[79] = t[108] ^ x[39];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[109] ^ x[43];
  assign t[81] = t[110] ^ x[45];
  assign t[82] = t[111] ^ x[47];
  assign t[83] = t[112] ^ x[49];
  assign t[84] = t[113] ^ x[51];
  assign t[85] = t[114] ^ x[54];
  assign t[86] = t[115] ^ x[56];
  assign t[87] = t[116] ^ x[58];
  assign t[88] = t[117] ^ x[61];
  assign t[89] = t[118] ^ x[63];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[119] ^ x[65];
  assign t[91] = t[120] ^ x[67];
  assign t[92] = t[121] ^ x[69];
  assign t[93] = t[122] ^ x[71];
  assign t[94] = t[123] ^ x[73];
  assign t[95] = t[124] ^ x[75];
  assign t[96] = t[125] ^ x[77];
  assign t[97] = t[126] ^ x[79];
  assign t[98] = (x[0] & x[1]);
  assign t[99] = (x[8] & x[9]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[69];
endmodule

module R1ind131(x, y);
 input [79:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[129] ^ x[73];
  assign t[101] = t[130] ^ x[75];
  assign t[102] = t[131] ^ x[77];
  assign t[103] = t[132] ^ x[79];
  assign t[104] = (x[0] & x[1]);
  assign t[105] = (x[8] & x[9]);
  assign t[106] = (x[11] & x[12]);
  assign t[107] = (x[14] & x[15]);
  assign t[108] = (x[17] & x[18]);
  assign t[109] = (x[20] & x[21]);
  assign t[10] = ~(x[3]);
  assign t[110] = (x[20] & x[25]);
  assign t[111] = (x[20] & x[27]);
  assign t[112] = (x[29] & x[30]);
  assign t[113] = (x[32] & x[33]);
  assign t[114] = (x[37] & x[38]);
  assign t[115] = (x[20] & x[42]);
  assign t[116] = (x[29] & x[44]);
  assign t[117] = (x[29] & x[46]);
  assign t[118] = (x[32] & x[48]);
  assign t[119] = (x[32] & x[50]);
  assign t[11] = t[16] ? x[7] : x[6];
  assign t[120] = (x[52] & x[53]);
  assign t[121] = (x[37] & x[55]);
  assign t[122] = (x[37] & x[57]);
  assign t[123] = (x[59] & x[60]);
  assign t[124] = (x[29] & x[62]);
  assign t[125] = (x[32] & x[64]);
  assign t[126] = (x[52] & x[66]);
  assign t[127] = (x[52] & x[68]);
  assign t[128] = (x[37] & x[70]);
  assign t[129] = (x[59] & x[72]);
  assign t[12] = x[4] ? t[18] : t[17];
  assign t[130] = (x[59] & x[74]);
  assign t[131] = (x[52] & x[76]);
  assign t[132] = (x[59] & x[78]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[14] = ~(t[76] & t[77]);
  assign t[15] = ~(t[78] & t[79]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = t[24] ^ t[25];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = x[4] ? t[29] : t[28];
  assign t[21] = ~(t[78]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = ~(t[32] & t[80]);
  assign t[24] = t[16] ? x[24] : x[23];
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = ~(t[35] & t[36]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[81]);
  assign t[31] = ~(t[82]);
  assign t[32] = ~(t[43] & t[44]);
  assign t[33] = ~(t[45] & t[46]);
  assign t[34] = ~(t[47] & t[83]);
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = ~(t[50] & t[84]);
  assign t[37] = t[51] ? x[36] : x[35];
  assign t[38] = ~(t[52] & t[53]);
  assign t[39] = ~(t[54] & t[55]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[56] & t[85]);
  assign t[41] = t[16] ? x[41] : x[40];
  assign t[42] = ~(t[57] & t[58]);
  assign t[43] = ~(t[82] & t[81]);
  assign t[44] = ~(t[86]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[88]);
  assign t[47] = ~(t[59] & t[60]);
  assign t[48] = ~(t[89]);
  assign t[49] = ~(t[90]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[61] & t[62]);
  assign t[51] = ~(t[21]);
  assign t[52] = ~(t[63] & t[64]);
  assign t[53] = ~(t[65] & t[91]);
  assign t[54] = ~(t[92]);
  assign t[55] = ~(t[93]);
  assign t[56] = ~(t[66] & t[67]);
  assign t[57] = ~(t[68] & t[69]);
  assign t[58] = ~(t[70] & t[94]);
  assign t[59] = ~(t[88] & t[87]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95]);
  assign t[61] = ~(t[90] & t[89]);
  assign t[62] = ~(t[96]);
  assign t[63] = ~(t[97]);
  assign t[64] = ~(t[98]);
  assign t[65] = ~(t[71] & t[72]);
  assign t[66] = ~(t[93] & t[92]);
  assign t[67] = ~(t[99]);
  assign t[68] = ~(t[100]);
  assign t[69] = ~(t[101]);
  assign t[6] = t[11] ^ t[7];
  assign t[70] = ~(t[73] & t[74]);
  assign t[71] = ~(t[98] & t[97]);
  assign t[72] = ~(t[102]);
  assign t[73] = ~(t[101] & t[100]);
  assign t[74] = ~(t[103]);
  assign t[75] = t[104] ^ x[2];
  assign t[76] = t[105] ^ x[10];
  assign t[77] = t[106] ^ x[13];
  assign t[78] = t[107] ^ x[16];
  assign t[79] = t[108] ^ x[19];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[109] ^ x[22];
  assign t[81] = t[110] ^ x[26];
  assign t[82] = t[111] ^ x[28];
  assign t[83] = t[112] ^ x[31];
  assign t[84] = t[113] ^ x[34];
  assign t[85] = t[114] ^ x[39];
  assign t[86] = t[115] ^ x[43];
  assign t[87] = t[116] ^ x[45];
  assign t[88] = t[117] ^ x[47];
  assign t[89] = t[118] ^ x[49];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[119] ^ x[51];
  assign t[91] = t[120] ^ x[54];
  assign t[92] = t[121] ^ x[56];
  assign t[93] = t[122] ^ x[58];
  assign t[94] = t[123] ^ x[61];
  assign t[95] = t[124] ^ x[63];
  assign t[96] = t[125] ^ x[65];
  assign t[97] = t[126] ^ x[67];
  assign t[98] = t[127] ^ x[69];
  assign t[99] = t[128] ^ x[71];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[75];
endmodule

module R1ind132(x, y);
 input [67:0] x;
 output y;

 wire [108:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = (x[29] & x[48]);
  assign t[101] = (x[34] & x[50]);
  assign t[102] = (x[52] & x[53]);
  assign t[103] = (x[52] & x[55]);
  assign t[104] = (x[41] & x[57]);
  assign t[105] = (x[59] & x[60]);
  assign t[106] = (x[59] & x[62]);
  assign t[107] = (x[52] & x[64]);
  assign t[108] = (x[59] & x[66]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[7] : x[6];
  assign t[12] = x[4] ? t[18] : t[17];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[14] = ~(t[64] & t[65]);
  assign t[15] = ~(t[66] & t[67]);
  assign t[16] = ~(t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = t[24] ^ t[25];
  assign t[19] = x[4] ? t[27] : t[26];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = x[4] ? t[29] : t[28];
  assign t[21] = ~(t[66]);
  assign t[22] = ~(t[68] & t[30]);
  assign t[23] = ~(t[69] & t[31]);
  assign t[24] = t[16] ? x[26] : x[25];
  assign t[25] = ~(t[32] & t[33]);
  assign t[26] = ~(t[34] & t[35]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = ~(t[38] & t[39]);
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[70]);
  assign t[31] = ~(t[70] & t[42]);
  assign t[32] = ~(t[71] & t[43]);
  assign t[33] = ~(t[72] & t[44]);
  assign t[34] = ~(t[73] & t[45]);
  assign t[35] = ~(t[74] & t[46]);
  assign t[36] = t[47] ? x[40] : x[39];
  assign t[37] = ~(t[48] & t[49]);
  assign t[38] = ~(t[75] & t[50]);
  assign t[39] = ~(t[76] & t[51]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[16] ? x[47] : x[46];
  assign t[41] = ~(t[52] & t[53]);
  assign t[42] = ~(t[68]);
  assign t[43] = ~(t[77]);
  assign t[44] = ~(t[77] & t[54]);
  assign t[45] = ~(t[78]);
  assign t[46] = ~(t[78] & t[55]);
  assign t[47] = ~(t[21]);
  assign t[48] = ~(t[79] & t[56]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[81]);
  assign t[51] = ~(t[81] & t[58]);
  assign t[52] = ~(t[82] & t[59]);
  assign t[53] = ~(t[83] & t[60]);
  assign t[54] = ~(t[71]);
  assign t[55] = ~(t[73]);
  assign t[56] = ~(t[84]);
  assign t[57] = ~(t[84] & t[61]);
  assign t[58] = ~(t[75]);
  assign t[59] = ~(t[85]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[85] & t[62]);
  assign t[61] = ~(t[79]);
  assign t[62] = ~(t[82]);
  assign t[63] = t[86] ^ x[2];
  assign t[64] = t[87] ^ x[10];
  assign t[65] = t[88] ^ x[13];
  assign t[66] = t[89] ^ x[16];
  assign t[67] = t[90] ^ x[19];
  assign t[68] = t[91] ^ x[22];
  assign t[69] = t[92] ^ x[24];
  assign t[6] = t[11] ^ t[7];
  assign t[70] = t[93] ^ x[28];
  assign t[71] = t[94] ^ x[31];
  assign t[72] = t[95] ^ x[33];
  assign t[73] = t[96] ^ x[36];
  assign t[74] = t[97] ^ x[38];
  assign t[75] = t[98] ^ x[43];
  assign t[76] = t[99] ^ x[45];
  assign t[77] = t[100] ^ x[49];
  assign t[78] = t[101] ^ x[51];
  assign t[79] = t[102] ^ x[54];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[103] ^ x[56];
  assign t[81] = t[104] ^ x[58];
  assign t[82] = t[105] ^ x[61];
  assign t[83] = t[106] ^ x[63];
  assign t[84] = t[107] ^ x[65];
  assign t[85] = t[108] ^ x[67];
  assign t[86] = (x[0] & x[1]);
  assign t[87] = (x[8] & x[9]);
  assign t[88] = (x[11] & x[12]);
  assign t[89] = (x[14] & x[15]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = (x[17] & x[18]);
  assign t[91] = (x[20] & x[21]);
  assign t[92] = (x[20] & x[23]);
  assign t[93] = (x[20] & x[27]);
  assign t[94] = (x[29] & x[30]);
  assign t[95] = (x[29] & x[32]);
  assign t[96] = (x[34] & x[35]);
  assign t[97] = (x[34] & x[37]);
  assign t[98] = (x[41] & x[42]);
  assign t[99] = (x[41] & x[44]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[63];
endmodule

module R1ind133(x, y);
 input [79:0] x;
 output y;

 wire [201:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[161] | t[162]);
  assign t[101] = ~(t[169]);
  assign t[102] = ~(t[170]);
  assign t[103] = ~(t[124] | t[125]);
  assign t[104] = ~(t[33]);
  assign t[105] = ~(t[84] | t[126]);
  assign t[106] = ~(t[127]);
  assign t[107] = x[4] & t[146];
  assign t[108] = ~(t[148]);
  assign t[109] = ~(x[4] | t[146]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[146] | t[148]);
  assign t[111] = ~(x[4] | t[128]);
  assign t[112] = t[145] ? t[129] : t[83];
  assign t[113] = t[145] ? t[80] : t[130];
  assign t[114] = t[145] ? t[80] : t[81];
  assign t[115] = ~(t[34] | t[131]);
  assign t[116] = ~(t[53] & t[132]);
  assign t[117] = ~(t[122] & t[133]);
  assign t[118] = t[53] | t[134];
  assign t[119] = ~(t[171]);
  assign t[11] = ~(t[16] ^ t[17]);
  assign t[120] = ~(t[166] | t[167]);
  assign t[121] = ~(t[57] | t[135]);
  assign t[122] = t[148] & t[136];
  assign t[123] = ~(t[64]);
  assign t[124] = ~(t[172]);
  assign t[125] = ~(t[169] | t[170]);
  assign t[126] = ~(t[137] & t[64]);
  assign t[127] = ~(t[57] | t[138]);
  assign t[128] = ~(t[146]);
  assign t[129] = ~(x[4] & t[139]);
  assign t[12] = x[4] ? t[19] : t[18];
  assign t[130] = ~(t[109] & t[148]);
  assign t[131] = ~(t[57] | t[140]);
  assign t[132] = ~(t[82] & t[86]);
  assign t[133] = t[109] | t[107];
  assign t[134] = t[145] ? t[82] : t[83];
  assign t[135] = t[145] ? t[82] : t[86];
  assign t[136] = ~(t[53] | t[145]);
  assign t[137] = ~(t[141] | t[90]);
  assign t[138] = t[145] ? t[81] : t[142];
  assign t[139] = ~(t[146] | t[108]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[145] ? t[83] : t[129];
  assign t[141] = ~(t[57] | t[143]);
  assign t[142] = ~(t[107] & t[148]);
  assign t[143] = t[145] ? t[142] : t[81];
  assign t[144] = t[173] ^ x[2];
  assign t[145] = t[174] ^ x[10];
  assign t[146] = t[175] ^ x[13];
  assign t[147] = t[176] ^ x[16];
  assign t[148] = t[177] ^ x[19];
  assign t[149] = t[178] ^ x[22];
  assign t[14] = ~(t[145] & t[146]);
  assign t[150] = t[179] ^ x[24];
  assign t[151] = t[180] ^ x[26];
  assign t[152] = t[181] ^ x[29];
  assign t[153] = t[182] ^ x[34];
  assign t[154] = t[183] ^ x[37];
  assign t[155] = t[184] ^ x[39];
  assign t[156] = t[185] ^ x[41];
  assign t[157] = t[186] ^ x[43];
  assign t[158] = t[187] ^ x[45];
  assign t[159] = t[188] ^ x[47];
  assign t[15] = ~(t[147] & t[148]);
  assign t[160] = t[189] ^ x[50];
  assign t[161] = t[190] ^ x[54];
  assign t[162] = t[191] ^ x[56];
  assign t[163] = t[192] ^ x[59];
  assign t[164] = t[193] ^ x[63];
  assign t[165] = t[194] ^ x[65];
  assign t[166] = t[195] ^ x[67];
  assign t[167] = t[196] ^ x[69];
  assign t[168] = t[197] ^ x[71];
  assign t[169] = t[198] ^ x[73];
  assign t[16] = t[22] ? x[7] : x[6];
  assign t[170] = t[199] ^ x[75];
  assign t[171] = t[200] ^ x[77];
  assign t[172] = t[201] ^ x[79];
  assign t[173] = (x[0] & x[1]);
  assign t[174] = (x[8] & x[9]);
  assign t[175] = (x[11] & x[12]);
  assign t[176] = (x[14] & x[15]);
  assign t[177] = (x[17] & x[18]);
  assign t[178] = (x[20] & x[21]);
  assign t[179] = (x[20] & x[23]);
  assign t[17] = ~(t[23] & t[24]);
  assign t[180] = (x[20] & x[25]);
  assign t[181] = (x[27] & x[28]);
  assign t[182] = (x[32] & x[33]);
  assign t[183] = (x[35] & x[36]);
  assign t[184] = (x[20] & x[38]);
  assign t[185] = (x[27] & x[40]);
  assign t[186] = (x[27] & x[42]);
  assign t[187] = (x[32] & x[44]);
  assign t[188] = (x[32] & x[46]);
  assign t[189] = (x[48] & x[49]);
  assign t[18] = ~(t[25] | t[26]);
  assign t[190] = (x[35] & x[53]);
  assign t[191] = (x[35] & x[55]);
  assign t[192] = (x[57] & x[58]);
  assign t[193] = (x[27] & x[62]);
  assign t[194] = (x[32] & x[64]);
  assign t[195] = (x[48] & x[66]);
  assign t[196] = (x[48] & x[68]);
  assign t[197] = (x[35] & x[70]);
  assign t[198] = (x[57] & x[72]);
  assign t[199] = (x[57] & x[74]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[48] & x[76]);
  assign t[201] = (x[57] & x[78]);
  assign t[20] = x[4] ? t[30] : t[29];
  assign t[21] = x[4] ? t[32] : t[31];
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[34] | t[35]);
  assign t[24] = ~(t[36] | t[37]);
  assign t[25] = ~(t[38] | t[39]);
  assign t[26] = ~(t[149] | t[40]);
  assign t[27] = ~(t[41] | t[42]);
  assign t[28] = ~(t[43] ^ t[44]);
  assign t[29] = ~(t[45] | t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] ^ t[48]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[32] = ~(t[51] ^ t[52]);
  assign t[33] = ~(t[147]);
  assign t[34] = ~(t[53] | t[54]);
  assign t[35] = ~(t[53] | t[55]);
  assign t[36] = ~(t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = ~(t[150]);
  assign t[39] = ~(t[151]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] | t[60]);
  assign t[41] = ~(t[61] | t[62]);
  assign t[42] = ~(t[152] | t[63]);
  assign t[43] = t[22] ? x[31] : x[30];
  assign t[44] = ~(t[64] & t[65]);
  assign t[45] = ~(t[66] | t[67]);
  assign t[46] = ~(t[153] | t[68]);
  assign t[47] = ~(t[69] | t[70]);
  assign t[48] = ~(t[71] ^ t[72]);
  assign t[49] = ~(t[73] | t[74]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[154] | t[75]);
  assign t[51] = ~(t[76] | t[77]);
  assign t[52] = ~(t[78] ^ t[79]);
  assign t[53] = ~(t[147]);
  assign t[54] = t[145] ? t[81] : t[80];
  assign t[55] = t[145] ? t[83] : t[82];
  assign t[56] = ~(t[84] | t[85]);
  assign t[57] = ~(t[53]);
  assign t[58] = t[145] ? t[86] : t[82];
  assign t[59] = ~(t[155]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[150] | t[151]);
  assign t[61] = ~(t[156]);
  assign t[62] = ~(t[157]);
  assign t[63] = ~(t[87] | t[88]);
  assign t[64] = ~(t[89] | t[35]);
  assign t[65] = ~(t[90] | t[91]);
  assign t[66] = ~(t[158]);
  assign t[67] = ~(t[159]);
  assign t[68] = ~(t[92] | t[93]);
  assign t[69] = ~(t[94] | t[95]);
  assign t[6] = ~(t[7] ^ t[11]);
  assign t[70] = ~(t[160] | t[96]);
  assign t[71] = t[22] ? x[52] : x[51];
  assign t[72] = ~(t[97] & t[98]);
  assign t[73] = ~(t[161]);
  assign t[74] = ~(t[162]);
  assign t[75] = ~(t[99] | t[100]);
  assign t[76] = ~(t[101] | t[102]);
  assign t[77] = ~(t[163] | t[103]);
  assign t[78] = t[104] ? x[61] : x[60];
  assign t[79] = ~(t[105] & t[106]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[107] & t[108]);
  assign t[81] = ~(t[109] & t[108]);
  assign t[82] = ~(x[4] & t[110]);
  assign t[83] = ~(t[111] & t[108]);
  assign t[84] = ~(t[57] | t[112]);
  assign t[85] = ~(t[57] | t[113]);
  assign t[86] = ~(t[148] & t[111]);
  assign t[87] = ~(t[164]);
  assign t[88] = ~(t[156] | t[157]);
  assign t[89] = ~(t[53] | t[114]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[115] & t[116]);
  assign t[91] = ~(t[117] & t[118]);
  assign t[92] = ~(t[165]);
  assign t[93] = ~(t[158] | t[159]);
  assign t[94] = ~(t[166]);
  assign t[95] = ~(t[167]);
  assign t[96] = ~(t[119] | t[120]);
  assign t[97] = ~(t[121] | t[85]);
  assign t[98] = ~(t[122] | t[123]);
  assign t[99] = ~(t[168]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[144];
endmodule

module R1ind134(x, y);
 input [112:0] x;
 output y;

 wire [183:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = t[143] ^ x[2];
  assign t[103] = t[144] ^ x[10];
  assign t[104] = t[145] ^ x[13];
  assign t[105] = t[146] ^ x[16];
  assign t[106] = t[147] ^ x[19];
  assign t[107] = t[148] ^ x[22];
  assign t[108] = t[149] ^ x[27];
  assign t[109] = t[150] ^ x[31];
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[33];
  assign t[111] = t[152] ^ x[36];
  assign t[112] = t[153] ^ x[39];
  assign t[113] = t[154] ^ x[44];
  assign t[114] = t[155] ^ x[48];
  assign t[115] = t[156] ^ x[50];
  assign t[116] = t[157] ^ x[53];
  assign t[117] = t[158] ^ x[58];
  assign t[118] = t[159] ^ x[62];
  assign t[119] = t[160] ^ x[64];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[161] ^ x[66];
  assign t[121] = t[162] ^ x[68];
  assign t[122] = t[163] ^ x[70];
  assign t[123] = t[164] ^ x[72];
  assign t[124] = t[165] ^ x[74];
  assign t[125] = t[166] ^ x[76];
  assign t[126] = t[167] ^ x[78];
  assign t[127] = t[168] ^ x[80];
  assign t[128] = t[169] ^ x[83];
  assign t[129] = t[170] ^ x[85];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[87];
  assign t[131] = t[172] ^ x[90];
  assign t[132] = t[173] ^ x[92];
  assign t[133] = t[174] ^ x[94];
  assign t[134] = t[175] ^ x[96];
  assign t[135] = t[176] ^ x[98];
  assign t[136] = t[177] ^ x[100];
  assign t[137] = t[178] ^ x[102];
  assign t[138] = t[179] ^ x[104];
  assign t[139] = t[180] ^ x[106];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[108];
  assign t[141] = t[182] ^ x[110];
  assign t[142] = t[183] ^ x[112];
  assign t[143] = (x[0] & x[1]);
  assign t[144] = (x[8] & x[9]);
  assign t[145] = (x[11] & x[12]);
  assign t[146] = (x[14] & x[15]);
  assign t[147] = (x[17] & x[18]);
  assign t[148] = (x[20] & x[21]);
  assign t[149] = (x[25] & x[26]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[20] & x[30]);
  assign t[151] = (x[20] & x[32]);
  assign t[152] = (x[34] & x[35]);
  assign t[153] = (x[37] & x[38]);
  assign t[154] = (x[42] & x[43]);
  assign t[155] = (x[25] & x[47]);
  assign t[156] = (x[25] & x[49]);
  assign t[157] = (x[51] & x[52]);
  assign t[158] = (x[56] & x[57]);
  assign t[159] = (x[20] & x[61]);
  assign t[15] = ~(t[103] & t[104]);
  assign t[160] = (x[34] & x[63]);
  assign t[161] = (x[34] & x[65]);
  assign t[162] = (x[37] & x[67]);
  assign t[163] = (x[37] & x[69]);
  assign t[164] = (x[42] & x[71]);
  assign t[165] = (x[42] & x[73]);
  assign t[166] = (x[25] & x[75]);
  assign t[167] = (x[51] & x[77]);
  assign t[168] = (x[51] & x[79]);
  assign t[169] = (x[81] & x[82]);
  assign t[16] = ~(t[105] & t[106]);
  assign t[170] = (x[56] & x[84]);
  assign t[171] = (x[56] & x[86]);
  assign t[172] = (x[88] & x[89]);
  assign t[173] = (x[34] & x[91]);
  assign t[174] = (x[37] & x[93]);
  assign t[175] = (x[42] & x[95]);
  assign t[176] = (x[51] & x[97]);
  assign t[177] = (x[81] & x[99]);
  assign t[178] = (x[81] & x[101]);
  assign t[179] = (x[56] & x[103]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[88] & x[105]);
  assign t[181] = (x[88] & x[107]);
  assign t[182] = (x[81] & x[109]);
  assign t[183] = (x[88] & x[111]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[105]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[25];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] | t[107];
  assign t[31] = t[47] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[35];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[42];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = t[58] | t[108];
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = t[61] ^ t[62];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[109]);
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[67] | t[44]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[68] & t[69]);
  assign t[49] = t[70] | t[111];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[71] & t[72]);
  assign t[51] = t[73] | t[112];
  assign t[52] = t[74] ? x[41] : x[40];
  assign t[53] = ~(t[75] & t[76]);
  assign t[54] = t[77] | t[113];
  assign t[55] = t[74] ? x[46] : x[45];
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[78] | t[56]);
  assign t[59] = ~(t[79] & t[80]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[81] | t[116];
  assign t[61] = t[74] ? x[55] : x[54];
  assign t[62] = ~(t[82] & t[83]);
  assign t[63] = ~(t[84] & t[85]);
  assign t[64] = t[86] | t[117];
  assign t[65] = t[17] ? x[60] : x[59];
  assign t[66] = ~(t[87] & t[88]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[89] | t[68]);
  assign t[71] = ~(t[121]);
  assign t[72] = ~(t[122]);
  assign t[73] = ~(t[90] | t[71]);
  assign t[74] = ~(t[24]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[91] | t[75]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[92] | t[79]);
  assign t[82] = ~(t[93] & t[94]);
  assign t[83] = t[95] | t[128];
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[96] | t[84]);
  assign t[87] = ~(t[97] & t[98]);
  assign t[88] = t[99] | t[131];
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[136]);
  assign t[94] = ~(t[137]);
  assign t[95] = ~(t[100] | t[93]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[101] | t[97]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[102];
endmodule

module R1ind135(x, y);
 input [112:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[107] & t[108]);
  assign t[102] = ~(t[139] & t[138]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[109] & t[110]);
  assign t[107] = ~(t[146] & t[145]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[151]);
  assign t[111] = t[152] ^ x[2];
  assign t[112] = t[153] ^ x[10];
  assign t[113] = t[154] ^ x[13];
  assign t[114] = t[155] ^ x[16];
  assign t[115] = t[156] ^ x[19];
  assign t[116] = t[157] ^ x[22];
  assign t[117] = t[158] ^ x[27];
  assign t[118] = t[159] ^ x[31];
  assign t[119] = t[160] ^ x[33];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[161] ^ x[36];
  assign t[121] = t[162] ^ x[39];
  assign t[122] = t[163] ^ x[44];
  assign t[123] = t[164] ^ x[48];
  assign t[124] = t[165] ^ x[50];
  assign t[125] = t[166] ^ x[53];
  assign t[126] = t[167] ^ x[58];
  assign t[127] = t[168] ^ x[62];
  assign t[128] = t[169] ^ x[64];
  assign t[129] = t[170] ^ x[66];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[68];
  assign t[131] = t[172] ^ x[70];
  assign t[132] = t[173] ^ x[72];
  assign t[133] = t[174] ^ x[74];
  assign t[134] = t[175] ^ x[76];
  assign t[135] = t[176] ^ x[78];
  assign t[136] = t[177] ^ x[80];
  assign t[137] = t[178] ^ x[83];
  assign t[138] = t[179] ^ x[85];
  assign t[139] = t[180] ^ x[87];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[90];
  assign t[141] = t[182] ^ x[92];
  assign t[142] = t[183] ^ x[94];
  assign t[143] = t[184] ^ x[96];
  assign t[144] = t[185] ^ x[98];
  assign t[145] = t[186] ^ x[100];
  assign t[146] = t[187] ^ x[102];
  assign t[147] = t[188] ^ x[104];
  assign t[148] = t[189] ^ x[106];
  assign t[149] = t[190] ^ x[108];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[191] ^ x[110];
  assign t[151] = t[192] ^ x[112];
  assign t[152] = (x[0] & x[1]);
  assign t[153] = (x[8] & x[9]);
  assign t[154] = (x[11] & x[12]);
  assign t[155] = (x[14] & x[15]);
  assign t[156] = (x[17] & x[18]);
  assign t[157] = (x[20] & x[21]);
  assign t[158] = (x[25] & x[26]);
  assign t[159] = (x[20] & x[30]);
  assign t[15] = ~(t[112] & t[113]);
  assign t[160] = (x[20] & x[32]);
  assign t[161] = (x[34] & x[35]);
  assign t[162] = (x[37] & x[38]);
  assign t[163] = (x[42] & x[43]);
  assign t[164] = (x[25] & x[47]);
  assign t[165] = (x[25] & x[49]);
  assign t[166] = (x[51] & x[52]);
  assign t[167] = (x[56] & x[57]);
  assign t[168] = (x[20] & x[61]);
  assign t[169] = (x[34] & x[63]);
  assign t[16] = ~(t[114] & t[115]);
  assign t[170] = (x[34] & x[65]);
  assign t[171] = (x[37] & x[67]);
  assign t[172] = (x[37] & x[69]);
  assign t[173] = (x[42] & x[71]);
  assign t[174] = (x[42] & x[73]);
  assign t[175] = (x[25] & x[75]);
  assign t[176] = (x[51] & x[77]);
  assign t[177] = (x[51] & x[79]);
  assign t[178] = (x[81] & x[82]);
  assign t[179] = (x[56] & x[84]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[56] & x[86]);
  assign t[181] = (x[88] & x[89]);
  assign t[182] = (x[34] & x[91]);
  assign t[183] = (x[37] & x[93]);
  assign t[184] = (x[42] & x[95]);
  assign t[185] = (x[51] & x[97]);
  assign t[186] = (x[81] & x[99]);
  assign t[187] = (x[81] & x[101]);
  assign t[188] = (x[56] & x[103]);
  assign t[189] = (x[88] & x[105]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[88] & x[107]);
  assign t[191] = (x[81] & x[109]);
  assign t[192] = (x[88] & x[111]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[114]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[25];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[116]);
  assign t[31] = t[47] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[35];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[42];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = ~(t[58] & t[117]);
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = t[61] ^ t[62];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[118]);
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[67] & t[68]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = ~(t[71] & t[120]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = ~(t[74] & t[121]);
  assign t[52] = t[75] ? x[41] : x[40];
  assign t[53] = ~(t[76] & t[77]);
  assign t[54] = ~(t[78] & t[122]);
  assign t[55] = t[75] ? x[46] : x[45];
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[124]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[83] & t[125]);
  assign t[61] = t[75] ? x[55] : x[54];
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[88] & t[126]);
  assign t[65] = t[17] ? x[60] : x[59];
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = ~(t[119] & t[118]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[128]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[129]);
  assign t[71] = ~(t[91] & t[92]);
  assign t[72] = ~(t[130]);
  assign t[73] = ~(t[131]);
  assign t[74] = ~(t[93] & t[94]);
  assign t[75] = ~(t[24]);
  assign t[76] = ~(t[132]);
  assign t[77] = ~(t[133]);
  assign t[78] = ~(t[95] & t[96]);
  assign t[79] = ~(t[124] & t[123]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[97] & t[98]);
  assign t[84] = ~(t[99] & t[100]);
  assign t[85] = ~(t[101] & t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[102] & t[103]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[106] & t[140]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[131] & t[130]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[133] & t[132]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[136] & t[135]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[145]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[111];
endmodule

module R1ind136(x, y);
 input [94:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[29];
  assign t[101] = t[133] ^ x[31];
  assign t[102] = t[134] ^ x[35];
  assign t[103] = t[135] ^ x[38];
  assign t[104] = t[136] ^ x[40];
  assign t[105] = t[137] ^ x[43];
  assign t[106] = t[138] ^ x[45];
  assign t[107] = t[139] ^ x[50];
  assign t[108] = t[140] ^ x[52];
  assign t[109] = t[141] ^ x[56];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[59];
  assign t[111] = t[143] ^ x[61];
  assign t[112] = t[144] ^ x[66];
  assign t[113] = t[145] ^ x[68];
  assign t[114] = t[146] ^ x[72];
  assign t[115] = t[147] ^ x[74];
  assign t[116] = t[148] ^ x[76];
  assign t[117] = t[149] ^ x[78];
  assign t[118] = t[150] ^ x[81];
  assign t[119] = t[151] ^ x[83];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[152] ^ x[85];
  assign t[121] = t[153] ^ x[88];
  assign t[122] = t[154] ^ x[90];
  assign t[123] = t[155] ^ x[92];
  assign t[124] = t[156] ^ x[94];
  assign t[125] = (x[0] & x[1]);
  assign t[126] = (x[8] & x[9]);
  assign t[127] = (x[11] & x[12]);
  assign t[128] = (x[14] & x[15]);
  assign t[129] = (x[17] & x[18]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & x[21]);
  assign t[131] = (x[20] & x[23]);
  assign t[132] = (x[27] & x[28]);
  assign t[133] = (x[27] & x[30]);
  assign t[134] = (x[20] & x[34]);
  assign t[135] = (x[36] & x[37]);
  assign t[136] = (x[36] & x[39]);
  assign t[137] = (x[41] & x[42]);
  assign t[138] = (x[41] & x[44]);
  assign t[139] = (x[48] & x[49]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[48] & x[51]);
  assign t[141] = (x[27] & x[55]);
  assign t[142] = (x[57] & x[58]);
  assign t[143] = (x[57] & x[60]);
  assign t[144] = (x[64] & x[65]);
  assign t[145] = (x[64] & x[67]);
  assign t[146] = (x[36] & x[71]);
  assign t[147] = (x[41] & x[73]);
  assign t[148] = (x[48] & x[75]);
  assign t[149] = (x[57] & x[77]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[79] & x[80]);
  assign t[151] = (x[79] & x[82]);
  assign t[152] = (x[64] & x[84]);
  assign t[153] = (x[86] & x[87]);
  assign t[154] = (x[86] & x[89]);
  assign t[155] = (x[79] & x[91]);
  assign t[156] = (x[86] & x[93]);
  assign t[15] = ~(t[94] & t[95]);
  assign t[16] = ~(t[96] & t[97]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[96]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[25];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[98] & t[44]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = t[46] ? x[26] : x[25];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = t[51] ^ t[42];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[33];
  assign t[37] = ~(t[100] & t[55]);
  assign t[38] = ~(t[101] & t[56]);
  assign t[39] = t[17] ? x[33] : x[32];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = t[59] ^ t[60];
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[64];
  assign t[44] = ~(t[102]);
  assign t[45] = ~(t[102] & t[65]);
  assign t[46] = ~(t[24]);
  assign t[47] = ~(t[103] & t[66]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = ~(t[105] & t[68]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[106] & t[69]);
  assign t[51] = t[70] ? x[47] : x[46];
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = t[70] ? x[54] : x[53];
  assign t[55] = ~(t[109]);
  assign t[56] = ~(t[109] & t[73]);
  assign t[57] = ~(t[110] & t[74]);
  assign t[58] = ~(t[111] & t[75]);
  assign t[59] = t[70] ? x[63] : x[62];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[76] & t[77]);
  assign t[61] = ~(t[112] & t[78]);
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = t[17] ? x[70] : x[69];
  assign t[64] = ~(t[80] & t[81]);
  assign t[65] = ~(t[98]);
  assign t[66] = ~(t[114]);
  assign t[67] = ~(t[114] & t[82]);
  assign t[68] = ~(t[115]);
  assign t[69] = ~(t[115] & t[83]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[24]);
  assign t[71] = ~(t[116]);
  assign t[72] = ~(t[116] & t[84]);
  assign t[73] = ~(t[100]);
  assign t[74] = ~(t[117]);
  assign t[75] = ~(t[117] & t[85]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[107]);
  assign t[85] = ~(t[110]);
  assign t[86] = ~(t[123]);
  assign t[87] = ~(t[123] & t[91]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[124]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[124] & t[92]);
  assign t[91] = ~(t[118]);
  assign t[92] = ~(t[121]);
  assign t[93] = t[125] ^ x[2];
  assign t[94] = t[126] ^ x[10];
  assign t[95] = t[127] ^ x[13];
  assign t[96] = t[128] ^ x[16];
  assign t[97] = t[129] ^ x[19];
  assign t[98] = t[130] ^ x[22];
  assign t[99] = t[131] ^ x[24];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[93];
endmodule

module R1ind137(x, y);
 input [112:0] x;
 output y;

 wire [278:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[136] ? x[70] : x[69];
  assign t[101] = ~(t[141] & t[105]);
  assign t[102] = ~(t[220]);
  assign t[103] = ~(t[209] | t[210]);
  assign t[104] = ~(t[124] | t[49]);
  assign t[105] = ~(t[142] | t[138]);
  assign t[106] = ~(t[221]);
  assign t[107] = ~(t[222]);
  assign t[108] = ~(t[143] | t[144]);
  assign t[109] = ~(t[145] | t[146]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[223] | t[147]);
  assign t[111] = t[29] ? x[81] : x[80];
  assign t[112] = ~(t[148] & t[149]);
  assign t[113] = ~(t[224]);
  assign t[114] = ~(t[225]);
  assign t[115] = ~(t[150] | t[151]);
  assign t[116] = ~(t[152] | t[153]);
  assign t[117] = ~(t[226] | t[154]);
  assign t[118] = t[136] ? x[90] : x[89];
  assign t[119] = ~(t[155] & t[156]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[157] & t[158]);
  assign t[121] = ~(t[159] & t[158]);
  assign t[122] = ~(x[4] & t[160]);
  assign t[123] = ~(t[161] & t[158]);
  assign t[124] = ~(t[78] | t[162]);
  assign t[125] = ~(t[163] | t[164]);
  assign t[126] = ~(t[122] & t[165]);
  assign t[127] = t[201] & t[166];
  assign t[128] = t[157] | t[159];
  assign t[129] = t[198] ? t[122] : t[123];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[227]);
  assign t[131] = ~(t[214] | t[215]);
  assign t[132] = ~(t[167] & t[168]);
  assign t[133] = t[138] | t[169];
  assign t[134] = ~(t[228]);
  assign t[135] = ~(t[216] | t[217]);
  assign t[136] = ~(t[47]);
  assign t[137] = ~(t[30] & t[168]);
  assign t[138] = ~(t[163] | t[170]);
  assign t[139] = ~(t[229]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[218] | t[219]);
  assign t[141] = ~(t[171]);
  assign t[142] = ~(t[172]);
  assign t[143] = ~(t[230]);
  assign t[144] = ~(t[221] | t[222]);
  assign t[145] = ~(t[231]);
  assign t[146] = ~(t[232]);
  assign t[147] = ~(t[173] | t[174]);
  assign t[148] = ~(t[175] | t[176]);
  assign t[149] = ~(t[127] | t[177]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[233]);
  assign t[151] = ~(t[224] | t[225]);
  assign t[152] = ~(t[234]);
  assign t[153] = ~(t[235]);
  assign t[154] = ~(t[178] | t[179]);
  assign t[155] = ~(t[180] | t[181]);
  assign t[156] = ~(t[182]);
  assign t[157] = ~(x[4] | t[199]);
  assign t[158] = ~(t[201]);
  assign t[159] = x[4] & t[199];
  assign t[15] = ~(t[198] & t[199]);
  assign t[160] = ~(t[199] | t[201]);
  assign t[161] = ~(x[4] | t[183]);
  assign t[162] = t[198] ? t[120] : t[121];
  assign t[163] = ~(t[78]);
  assign t[164] = t[198] ? t[123] : t[184];
  assign t[165] = ~(t[201] & t[161]);
  assign t[166] = ~(t[78] | t[198]);
  assign t[167] = ~(t[166] & t[185]);
  assign t[168] = ~(t[186] & t[187]);
  assign t[169] = ~(t[163] | t[188]);
  assign t[16] = ~(t[200] & t[201]);
  assign t[170] = t[198] ? t[165] : t[122];
  assign t[171] = ~(t[163] | t[189]);
  assign t[172] = ~(t[180] | t[176]);
  assign t[173] = ~(t[236]);
  assign t[174] = ~(t[231] | t[232]);
  assign t[175] = ~(t[163] | t[190]);
  assign t[176] = ~(t[163] | t[191]);
  assign t[177] = ~(t[30]);
  assign t[178] = ~(t[237]);
  assign t[179] = ~(t[234] | t[235]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[163] | t[192]);
  assign t[181] = ~(t[193] & t[30]);
  assign t[182] = ~(t[163] | t[194]);
  assign t[183] = ~(t[199]);
  assign t[184] = ~(x[4] & t[186]);
  assign t[185] = ~(t[165] & t[184]);
  assign t[186] = ~(t[199] | t[158]);
  assign t[187] = t[163] & t[198];
  assign t[188] = t[198] ? t[195] : t[121];
  assign t[189] = t[198] ? t[196] : t[120];
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[198] ? t[122] : t[165];
  assign t[191] = t[198] ? t[121] : t[195];
  assign t[192] = t[198] ? t[184] : t[123];
  assign t[193] = ~(t[171] | t[50]);
  assign t[194] = t[198] ? t[120] : t[196];
  assign t[195] = ~(t[157] & t[201]);
  assign t[196] = ~(t[159] & t[201]);
  assign t[197] = t[238] ^ x[2];
  assign t[198] = t[239] ^ x[10];
  assign t[199] = t[240] ^ x[13];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[241] ^ x[16];
  assign t[201] = t[242] ^ x[19];
  assign t[202] = t[243] ^ x[22];
  assign t[203] = t[244] ^ x[25];
  assign t[204] = t[245] ^ x[27];
  assign t[205] = t[246] ^ x[29];
  assign t[206] = t[247] ^ x[32];
  assign t[207] = t[248] ^ x[37];
  assign t[208] = t[249] ^ x[40];
  assign t[209] = t[250] ^ x[42];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[251] ^ x[44];
  assign t[211] = t[252] ^ x[49];
  assign t[212] = t[253] ^ x[52];
  assign t[213] = t[254] ^ x[54];
  assign t[214] = t[255] ^ x[56];
  assign t[215] = t[256] ^ x[58];
  assign t[216] = t[257] ^ x[60];
  assign t[217] = t[258] ^ x[62];
  assign t[218] = t[259] ^ x[66];
  assign t[219] = t[260] ^ x[68];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[261] ^ x[72];
  assign t[221] = t[262] ^ x[74];
  assign t[222] = t[263] ^ x[76];
  assign t[223] = t[264] ^ x[79];
  assign t[224] = t[265] ^ x[83];
  assign t[225] = t[266] ^ x[85];
  assign t[226] = t[267] ^ x[88];
  assign t[227] = t[268] ^ x[92];
  assign t[228] = t[269] ^ x[94];
  assign t[229] = t[270] ^ x[96];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[271] ^ x[98];
  assign t[231] = t[272] ^ x[100];
  assign t[232] = t[273] ^ x[102];
  assign t[233] = t[274] ^ x[104];
  assign t[234] = t[275] ^ x[106];
  assign t[235] = t[276] ^ x[108];
  assign t[236] = t[277] ^ x[110];
  assign t[237] = t[278] ^ x[112];
  assign t[238] = (x[0] & x[1]);
  assign t[239] = (x[8] & x[9]);
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = (x[11] & x[12]);
  assign t[241] = (x[14] & x[15]);
  assign t[242] = (x[17] & x[18]);
  assign t[243] = (x[20] & x[21]);
  assign t[244] = (x[23] & x[24]);
  assign t[245] = (x[20] & x[26]);
  assign t[246] = (x[20] & x[28]);
  assign t[247] = (x[30] & x[31]);
  assign t[248] = (x[35] & x[36]);
  assign t[249] = (x[38] & x[39]);
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = (x[23] & x[41]);
  assign t[251] = (x[23] & x[43]);
  assign t[252] = (x[47] & x[48]);
  assign t[253] = (x[50] & x[51]);
  assign t[254] = (x[20] & x[53]);
  assign t[255] = (x[30] & x[55]);
  assign t[256] = (x[30] & x[57]);
  assign t[257] = (x[35] & x[59]);
  assign t[258] = (x[35] & x[61]);
  assign t[259] = (x[38] & x[65]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[38] & x[67]);
  assign t[261] = (x[23] & x[71]);
  assign t[262] = (x[47] & x[73]);
  assign t[263] = (x[47] & x[75]);
  assign t[264] = (x[77] & x[78]);
  assign t[265] = (x[50] & x[82]);
  assign t[266] = (x[50] & x[84]);
  assign t[267] = (x[86] & x[87]);
  assign t[268] = (x[30] & x[91]);
  assign t[269] = (x[35] & x[93]);
  assign t[26] = ~(t[25] ^ t[42]);
  assign t[270] = (x[38] & x[95]);
  assign t[271] = (x[47] & x[97]);
  assign t[272] = (x[77] & x[99]);
  assign t[273] = (x[77] & x[101]);
  assign t[274] = (x[50] & x[103]);
  assign t[275] = (x[86] & x[105]);
  assign t[276] = (x[86] & x[107]);
  assign t[277] = (x[77] & x[109]);
  assign t[278] = (x[86] & x[111]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[29] = ~(t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[202] | t[54]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[36] = ~(t[59] | t[60]);
  assign t[37] = ~(t[38] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[43] ^ t[64]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[65] | t[66]);
  assign t[41] = ~(t[203] | t[67]);
  assign t[42] = ~(t[68] ^ t[69]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[47] = ~(t[200]);
  assign t[48] = ~(t[78] | t[79]);
  assign t[49] = ~(t[78] | t[80]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[81] & t[82]);
  assign t[51] = ~(t[83] & t[84]);
  assign t[52] = ~(t[204]);
  assign t[53] = ~(t[205]);
  assign t[54] = ~(t[85] | t[86]);
  assign t[55] = ~(t[87] | t[88]);
  assign t[56] = ~(t[206] | t[89]);
  assign t[57] = t[90] ? x[34] : x[33];
  assign t[58] = ~(t[91] & t[83]);
  assign t[59] = ~(t[92] | t[93]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[207] | t[94]);
  assign t[61] = ~(t[95] ^ t[96]);
  assign t[62] = ~(t[97] | t[98]);
  assign t[63] = ~(t[208] | t[99]);
  assign t[64] = ~(t[100] ^ t[101]);
  assign t[65] = ~(t[209]);
  assign t[66] = ~(t[210]);
  assign t[67] = ~(t[102] | t[103]);
  assign t[68] = t[29] ? x[46] : x[45];
  assign t[69] = ~(t[104] & t[105]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[211] | t[108]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[111] ^ t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[212] | t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[200]);
  assign t[79] = t[198] ? t[121] : t[120];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[198] ? t[123] : t[122];
  assign t[81] = ~(t[124] | t[125]);
  assign t[82] = ~(t[78] & t[126]);
  assign t[83] = ~(t[127] & t[128]);
  assign t[84] = t[78] | t[129];
  assign t[85] = ~(t[213]);
  assign t[86] = ~(t[204] | t[205]);
  assign t[87] = ~(t[214]);
  assign t[88] = ~(t[215]);
  assign t[89] = ~(t[130] | t[131]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[47]);
  assign t[91] = ~(t[132] | t[133]);
  assign t[92] = ~(t[216]);
  assign t[93] = ~(t[217]);
  assign t[94] = ~(t[134] | t[135]);
  assign t[95] = t[136] ? x[64] : x[63];
  assign t[96] = t[137] | t[138];
  assign t[97] = ~(t[218]);
  assign t[98] = ~(t[219]);
  assign t[99] = ~(t[139] | t[140]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[197];
endmodule

module R1ind138(x, y);
 input [112:0] x;
 output y;

 wire [182:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141]);
  assign t[101] = t[142] ^ x[2];
  assign t[102] = t[143] ^ x[10];
  assign t[103] = t[144] ^ x[13];
  assign t[104] = t[145] ^ x[16];
  assign t[105] = t[146] ^ x[19];
  assign t[106] = t[147] ^ x[22];
  assign t[107] = t[148] ^ x[27];
  assign t[108] = t[149] ^ x[31];
  assign t[109] = t[150] ^ x[33];
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[36];
  assign t[111] = t[152] ^ x[41];
  assign t[112] = t[153] ^ x[45];
  assign t[113] = t[154] ^ x[47];
  assign t[114] = t[155] ^ x[50];
  assign t[115] = t[156] ^ x[53];
  assign t[116] = t[157] ^ x[58];
  assign t[117] = t[158] ^ x[62];
  assign t[118] = t[159] ^ x[64];
  assign t[119] = t[160] ^ x[66];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[161] ^ x[69];
  assign t[121] = t[162] ^ x[71];
  assign t[122] = t[163] ^ x[73];
  assign t[123] = t[164] ^ x[75];
  assign t[124] = t[165] ^ x[77];
  assign t[125] = t[166] ^ x[79];
  assign t[126] = t[167] ^ x[81];
  assign t[127] = t[168] ^ x[83];
  assign t[128] = t[169] ^ x[85];
  assign t[129] = t[170] ^ x[87];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[90];
  assign t[131] = t[172] ^ x[92];
  assign t[132] = t[173] ^ x[94];
  assign t[133] = t[174] ^ x[96];
  assign t[134] = t[175] ^ x[98];
  assign t[135] = t[176] ^ x[100];
  assign t[136] = t[177] ^ x[102];
  assign t[137] = t[178] ^ x[104];
  assign t[138] = t[179] ^ x[106];
  assign t[139] = t[180] ^ x[108];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[110];
  assign t[141] = t[182] ^ x[112];
  assign t[142] = (x[0] & x[1]);
  assign t[143] = (x[8] & x[9]);
  assign t[144] = (x[11] & x[12]);
  assign t[145] = (x[14] & x[15]);
  assign t[146] = (x[17] & x[18]);
  assign t[147] = (x[20] & x[21]);
  assign t[148] = (x[25] & x[26]);
  assign t[149] = (x[20] & x[30]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[20] & x[32]);
  assign t[151] = (x[34] & x[35]);
  assign t[152] = (x[39] & x[40]);
  assign t[153] = (x[25] & x[44]);
  assign t[154] = (x[25] & x[46]);
  assign t[155] = (x[48] & x[49]);
  assign t[156] = (x[51] & x[52]);
  assign t[157] = (x[56] & x[57]);
  assign t[158] = (x[20] & x[61]);
  assign t[159] = (x[34] & x[63]);
  assign t[15] = ~(t[102] & t[103]);
  assign t[160] = (x[34] & x[65]);
  assign t[161] = (x[67] & x[68]);
  assign t[162] = (x[39] & x[70]);
  assign t[163] = (x[39] & x[72]);
  assign t[164] = (x[25] & x[74]);
  assign t[165] = (x[48] & x[76]);
  assign t[166] = (x[48] & x[78]);
  assign t[167] = (x[51] & x[80]);
  assign t[168] = (x[51] & x[82]);
  assign t[169] = (x[56] & x[84]);
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = (x[56] & x[86]);
  assign t[171] = (x[88] & x[89]);
  assign t[172] = (x[34] & x[91]);
  assign t[173] = (x[67] & x[93]);
  assign t[174] = (x[67] & x[95]);
  assign t[175] = (x[39] & x[97]);
  assign t[176] = (x[48] & x[99]);
  assign t[177] = (x[51] & x[101]);
  assign t[178] = (x[56] & x[103]);
  assign t[179] = (x[88] & x[105]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[88] & x[107]);
  assign t[181] = (x[67] & x[109]);
  assign t[182] = (x[88] & x[111]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[25];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[104]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] | t[106];
  assign t[31] = t[104] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[50];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] | t[107];
  assign t[38] = t[57] ? x[29] : x[28];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[40];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[108]);
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[67] | t[44]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = t[70] | t[110];
  assign t[49] = t[104] ? x[38] : x[37];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[71] & t[72]);
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = t[75] | t[111];
  assign t[53] = t[104] ? x[43] : x[42];
  assign t[54] = ~(t[112]);
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[76] | t[54]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[77] & t[78]);
  assign t[59] = t[79] | t[114];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[80] & t[81]);
  assign t[61] = t[82] | t[115];
  assign t[62] = t[17] ? x[55] : x[54];
  assign t[63] = ~(t[83] & t[84]);
  assign t[64] = t[85] | t[116];
  assign t[65] = t[17] ? x[60] : x[59];
  assign t[66] = ~(t[86] & t[87]);
  assign t[67] = ~(t[117]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[119]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[88] | t[68]);
  assign t[71] = ~(t[89] & t[90]);
  assign t[72] = t[91] | t[120];
  assign t[73] = ~(t[121]);
  assign t[74] = ~(t[122]);
  assign t[75] = ~(t[92] | t[73]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[93] | t[77]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[94] | t[80]);
  assign t[83] = ~(t[128]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[95] | t[83]);
  assign t[86] = ~(t[96] & t[97]);
  assign t[87] = t[98] | t[130];
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[99] | t[89]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[100] | t[96]);
  assign t[99] = ~(t[140]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[101];
endmodule

module R1ind139(x, y);
 input [112:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[145]);
  assign t[101] = ~(t[138] & t[137]);
  assign t[102] = ~(t[146]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[108] & t[109]);
  assign t[106] = ~(t[142] & t[141]);
  assign t[107] = ~(t[149]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[150]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[2];
  assign t[111] = t[152] ^ x[10];
  assign t[112] = t[153] ^ x[13];
  assign t[113] = t[154] ^ x[16];
  assign t[114] = t[155] ^ x[19];
  assign t[115] = t[156] ^ x[22];
  assign t[116] = t[157] ^ x[27];
  assign t[117] = t[158] ^ x[31];
  assign t[118] = t[159] ^ x[33];
  assign t[119] = t[160] ^ x[36];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[161] ^ x[41];
  assign t[121] = t[162] ^ x[45];
  assign t[122] = t[163] ^ x[47];
  assign t[123] = t[164] ^ x[50];
  assign t[124] = t[165] ^ x[53];
  assign t[125] = t[166] ^ x[58];
  assign t[126] = t[167] ^ x[62];
  assign t[127] = t[168] ^ x[64];
  assign t[128] = t[169] ^ x[66];
  assign t[129] = t[170] ^ x[69];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[71];
  assign t[131] = t[172] ^ x[73];
  assign t[132] = t[173] ^ x[75];
  assign t[133] = t[174] ^ x[77];
  assign t[134] = t[175] ^ x[79];
  assign t[135] = t[176] ^ x[81];
  assign t[136] = t[177] ^ x[83];
  assign t[137] = t[178] ^ x[85];
  assign t[138] = t[179] ^ x[87];
  assign t[139] = t[180] ^ x[90];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[92];
  assign t[141] = t[182] ^ x[94];
  assign t[142] = t[183] ^ x[96];
  assign t[143] = t[184] ^ x[98];
  assign t[144] = t[185] ^ x[100];
  assign t[145] = t[186] ^ x[102];
  assign t[146] = t[187] ^ x[104];
  assign t[147] = t[188] ^ x[106];
  assign t[148] = t[189] ^ x[108];
  assign t[149] = t[190] ^ x[110];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[191] ^ x[112];
  assign t[151] = (x[0] & x[1]);
  assign t[152] = (x[8] & x[9]);
  assign t[153] = (x[11] & x[12]);
  assign t[154] = (x[14] & x[15]);
  assign t[155] = (x[17] & x[18]);
  assign t[156] = (x[20] & x[21]);
  assign t[157] = (x[25] & x[26]);
  assign t[158] = (x[20] & x[30]);
  assign t[159] = (x[20] & x[32]);
  assign t[15] = ~(t[111] & t[112]);
  assign t[160] = (x[34] & x[35]);
  assign t[161] = (x[39] & x[40]);
  assign t[162] = (x[25] & x[44]);
  assign t[163] = (x[25] & x[46]);
  assign t[164] = (x[48] & x[49]);
  assign t[165] = (x[51] & x[52]);
  assign t[166] = (x[56] & x[57]);
  assign t[167] = (x[20] & x[61]);
  assign t[168] = (x[34] & x[63]);
  assign t[169] = (x[34] & x[65]);
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = (x[67] & x[68]);
  assign t[171] = (x[39] & x[70]);
  assign t[172] = (x[39] & x[72]);
  assign t[173] = (x[25] & x[74]);
  assign t[174] = (x[48] & x[76]);
  assign t[175] = (x[48] & x[78]);
  assign t[176] = (x[51] & x[80]);
  assign t[177] = (x[51] & x[82]);
  assign t[178] = (x[56] & x[84]);
  assign t[179] = (x[56] & x[86]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[88] & x[89]);
  assign t[181] = (x[34] & x[91]);
  assign t[182] = (x[67] & x[93]);
  assign t[183] = (x[67] & x[95]);
  assign t[184] = (x[39] & x[97]);
  assign t[185] = (x[48] & x[99]);
  assign t[186] = (x[51] & x[101]);
  assign t[187] = (x[56] & x[103]);
  assign t[188] = (x[88] & x[105]);
  assign t[189] = (x[88] & x[107]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[67] & x[109]);
  assign t[191] = (x[88] & x[111]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[25];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[113]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[115]);
  assign t[31] = t[113] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[50];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = ~(t[56] & t[116]);
  assign t[38] = t[57] ? x[29] : x[28];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[40];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[117]);
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[67] & t[68]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = ~(t[71] & t[119]);
  assign t[49] = t[113] ? x[38] : x[37];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = ~(t[76] & t[120]);
  assign t[53] = t[113] ? x[43] : x[42];
  assign t[54] = ~(t[121]);
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[77] & t[78]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[81] & t[123]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = ~(t[84] & t[124]);
  assign t[62] = t[17] ? x[55] : x[54];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = ~(t[87] & t[125]);
  assign t[65] = t[17] ? x[60] : x[59];
  assign t[66] = ~(t[88] & t[89]);
  assign t[67] = ~(t[118] & t[117]);
  assign t[68] = ~(t[126]);
  assign t[69] = ~(t[127]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[90] & t[91]);
  assign t[72] = ~(t[92] & t[93]);
  assign t[73] = ~(t[94] & t[129]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[131]);
  assign t[76] = ~(t[95] & t[96]);
  assign t[77] = ~(t[122] & t[121]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[97] & t[98]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] & t[100]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[101] & t[102]);
  assign t[88] = ~(t[103] & t[104]);
  assign t[89] = ~(t[105] & t[139]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[106] & t[107]);
  assign t[95] = ~(t[131] & t[130]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[134] & t[133]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[110];
endmodule

module R1ind140(x, y);
 input [94:0] x;
 output y;

 wire [155:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[31];
  assign t[101] = t[133] ^ x[35];
  assign t[102] = t[134] ^ x[38];
  assign t[103] = t[135] ^ x[40];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[47];
  assign t[106] = t[138] ^ x[51];
  assign t[107] = t[139] ^ x[54];
  assign t[108] = t[140] ^ x[56];
  assign t[109] = t[141] ^ x[59];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[61];
  assign t[111] = t[143] ^ x[66];
  assign t[112] = t[144] ^ x[68];
  assign t[113] = t[145] ^ x[72];
  assign t[114] = t[146] ^ x[74];
  assign t[115] = t[147] ^ x[77];
  assign t[116] = t[148] ^ x[79];
  assign t[117] = t[149] ^ x[81];
  assign t[118] = t[150] ^ x[83];
  assign t[119] = t[151] ^ x[86];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[152] ^ x[88];
  assign t[121] = t[153] ^ x[90];
  assign t[122] = t[154] ^ x[92];
  assign t[123] = t[155] ^ x[94];
  assign t[124] = (x[0] & x[1]);
  assign t[125] = (x[8] & x[9]);
  assign t[126] = (x[11] & x[12]);
  assign t[127] = (x[14] & x[15]);
  assign t[128] = (x[17] & x[18]);
  assign t[129] = (x[20] & x[21]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & x[23]);
  assign t[131] = (x[27] & x[28]);
  assign t[132] = (x[27] & x[30]);
  assign t[133] = (x[20] & x[34]);
  assign t[134] = (x[36] & x[37]);
  assign t[135] = (x[36] & x[39]);
  assign t[136] = (x[43] & x[44]);
  assign t[137] = (x[43] & x[46]);
  assign t[138] = (x[27] & x[50]);
  assign t[139] = (x[52] & x[53]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[52] & x[55]);
  assign t[141] = (x[57] & x[58]);
  assign t[142] = (x[57] & x[60]);
  assign t[143] = (x[64] & x[65]);
  assign t[144] = (x[64] & x[67]);
  assign t[145] = (x[36] & x[71]);
  assign t[146] = (x[43] & x[73]);
  assign t[147] = (x[75] & x[76]);
  assign t[148] = (x[75] & x[78]);
  assign t[149] = (x[52] & x[80]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[57] & x[82]);
  assign t[151] = (x[84] & x[85]);
  assign t[152] = (x[84] & x[87]);
  assign t[153] = (x[64] & x[89]);
  assign t[154] = (x[75] & x[91]);
  assign t[155] = (x[84] & x[93]);
  assign t[15] = ~(t[93] & t[94]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[25];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[95]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[97] & t[44]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[98] & t[45]);
  assign t[31] = t[95] ? x[26] : x[25];
  assign t[32] = ~(t[46] & t[47]);
  assign t[33] = t[48] ^ t[32];
  assign t[34] = ~(t[49] & t[50]);
  assign t[35] = t[51] ^ t[52];
  assign t[36] = ~(t[99] & t[53]);
  assign t[37] = ~(t[100] & t[54]);
  assign t[38] = t[55] ? x[33] : x[32];
  assign t[39] = ~(t[56] & t[57]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = t[60] ^ t[61];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[42];
  assign t[44] = ~(t[101]);
  assign t[45] = ~(t[101] & t[65]);
  assign t[46] = ~(t[102] & t[66]);
  assign t[47] = ~(t[103] & t[67]);
  assign t[48] = t[95] ? x[42] : x[41];
  assign t[49] = ~(t[104] & t[68]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = t[95] ? x[49] : x[48];
  assign t[52] = ~(t[70] & t[71]);
  assign t[53] = ~(t[106]);
  assign t[54] = ~(t[106] & t[72]);
  assign t[55] = ~(t[24]);
  assign t[56] = ~(t[107] & t[73]);
  assign t[57] = ~(t[108] & t[74]);
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = ~(t[110] & t[76]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[17] ? x[63] : x[62];
  assign t[61] = ~(t[77] & t[78]);
  assign t[62] = ~(t[111] & t[79]);
  assign t[63] = ~(t[112] & t[80]);
  assign t[64] = t[17] ? x[70] : x[69];
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[113]);
  assign t[67] = ~(t[113] & t[81]);
  assign t[68] = ~(t[114]);
  assign t[69] = ~(t[114] & t[82]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[99]);
  assign t[73] = ~(t[117]);
  assign t[74] = ~(t[117] & t[85]);
  assign t[75] = ~(t[118]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[102]);
  assign t[82] = ~(t[104]);
  assign t[83] = ~(t[122]);
  assign t[84] = ~(t[122] & t[90]);
  assign t[85] = ~(t[107]);
  assign t[86] = ~(t[109]);
  assign t[87] = ~(t[123]);
  assign t[88] = ~(t[123] & t[91]);
  assign t[89] = ~(t[111]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[115]);
  assign t[91] = ~(t[119]);
  assign t[92] = t[124] ^ x[2];
  assign t[93] = t[125] ^ x[10];
  assign t[94] = t[126] ^ x[13];
  assign t[95] = t[127] ^ x[16];
  assign t[96] = t[128] ^ x[19];
  assign t[97] = t[129] ^ x[22];
  assign t[98] = t[130] ^ x[24];
  assign t[99] = t[131] ^ x[29];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[92];
endmodule

module R1ind141(x, y);
 input [112:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[211] | t[212]);
  assign t[101] = ~(t[223]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[139] | t[140]);
  assign t[104] = ~(t[47]);
  assign t[105] = ~(t[128] | t[141]);
  assign t[106] = ~(t[126]);
  assign t[107] = ~(t[225]);
  assign t[108] = ~(t[226]);
  assign t[109] = ~(t[142] | t[143]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[29] ? x[81] : x[80];
  assign t[111] = ~(t[144] & t[145]);
  assign t[112] = ~(t[227]);
  assign t[113] = ~(t[228]);
  assign t[114] = ~(t[146] | t[147]);
  assign t[115] = ~(t[148] | t[149]);
  assign t[116] = ~(t[229] | t[150]);
  assign t[117] = t[29] ? x[90] : x[89];
  assign t[118] = ~(t[82] & t[151]);
  assign t[119] = ~(t[203]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[204] & t[152]);
  assign t[121] = ~(x[4] & t[153]);
  assign t[122] = ~(t[154] & t[204]);
  assign t[123] = ~(t[155] & t[156]);
  assign t[124] = ~(t[119] | t[157]);
  assign t[125] = ~(t[119] | t[158]);
  assign t[126] = ~(t[78] | t[159]);
  assign t[127] = ~(t[160] & t[161]);
  assign t[128] = ~(t[78] | t[162]);
  assign t[129] = ~(t[230]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[217] | t[218]);
  assign t[131] = ~(t[231]);
  assign t[132] = ~(t[232]);
  assign t[133] = ~(t[163] | t[164]);
  assign t[134] = ~(t[137] | t[165]);
  assign t[135] = ~(t[233]);
  assign t[136] = ~(t[220] | t[221]);
  assign t[137] = ~(t[166] & t[167]);
  assign t[138] = ~(t[168] & t[30]);
  assign t[139] = ~(t[234]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[223] | t[224]);
  assign t[141] = ~(t[169] & t[82]);
  assign t[142] = ~(t[235]);
  assign t[143] = ~(t[225] | t[226]);
  assign t[144] = ~(t[170] | t[125]);
  assign t[145] = ~(t[171] | t[172]);
  assign t[146] = ~(t[236]);
  assign t[147] = ~(t[227] | t[228]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[238]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[173] | t[174]);
  assign t[151] = ~(t[175] | t[176]);
  assign t[152] = ~(x[4] | t[177]);
  assign t[153] = ~(t[202] | t[204]);
  assign t[154] = ~(x[4] | t[202]);
  assign t[155] = x[4] & t[202];
  assign t[156] = ~(t[204]);
  assign t[157] = t[201] ? t[123] : t[178];
  assign t[158] = t[201] ? t[179] : t[121];
  assign t[159] = t[201] ? t[178] : t[180];
  assign t[15] = ~(t[201] & t[202]);
  assign t[160] = ~(t[181] | t[48]);
  assign t[161] = ~(t[50] & t[182]);
  assign t[162] = t[201] ? t[183] : t[179];
  assign t[163] = ~(t[239]);
  assign t[164] = ~(t[231] | t[232]);
  assign t[165] = ~(t[184] & t[185]);
  assign t[166] = ~(t[81] & t[186]);
  assign t[167] = ~(t[187] & t[188]);
  assign t[168] = ~(t[126] | t[189]);
  assign t[169] = ~(t[181] | t[175]);
  assign t[16] = ~(t[203] & t[204]);
  assign t[170] = ~(t[119] | t[190]);
  assign t[171] = ~(t[86]);
  assign t[172] = ~(t[78] | t[191]);
  assign t[173] = ~(t[240]);
  assign t[174] = ~(t[237] | t[238]);
  assign t[175] = ~(t[192] & t[193]);
  assign t[176] = ~(t[161] & t[185]);
  assign t[177] = ~(t[202]);
  assign t[178] = ~(t[154] & t[156]);
  assign t[179] = ~(t[152] & t[156]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[155] & t[204]);
  assign t[181] = ~(t[78] | t[194]);
  assign t[182] = t[154] | t[155];
  assign t[183] = ~(x[4] & t[187]);
  assign t[184] = ~(t[125]);
  assign t[185] = t[119] | t[195];
  assign t[186] = ~(t[120] & t[183]);
  assign t[187] = ~(t[202] | t[156]);
  assign t[188] = t[78] & t[201];
  assign t[189] = ~(t[78] | t[196]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[201] ? t[178] : t[123];
  assign t[191] = t[201] ? t[120] : t[121];
  assign t[192] = ~(t[170] | t[197]);
  assign t[193] = ~(t[119] & t[198]);
  assign t[194] = t[201] ? t[180] : t[178];
  assign t[195] = t[201] ? t[121] : t[179];
  assign t[196] = t[201] ? t[122] : t[123];
  assign t[197] = ~(t[78] | t[199]);
  assign t[198] = ~(t[121] & t[120]);
  assign t[199] = t[201] ? t[179] : t[183];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[241] ^ x[2];
  assign t[201] = t[242] ^ x[10];
  assign t[202] = t[243] ^ x[13];
  assign t[203] = t[244] ^ x[16];
  assign t[204] = t[245] ^ x[19];
  assign t[205] = t[246] ^ x[22];
  assign t[206] = t[247] ^ x[25];
  assign t[207] = t[248] ^ x[27];
  assign t[208] = t[249] ^ x[29];
  assign t[209] = t[250] ^ x[34];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[251] ^ x[37];
  assign t[211] = t[252] ^ x[39];
  assign t[212] = t[253] ^ x[41];
  assign t[213] = t[254] ^ x[44];
  assign t[214] = t[255] ^ x[49];
  assign t[215] = t[256] ^ x[52];
  assign t[216] = t[257] ^ x[54];
  assign t[217] = t[258] ^ x[56];
  assign t[218] = t[259] ^ x[58];
  assign t[219] = t[260] ^ x[61];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[261] ^ x[65];
  assign t[221] = t[262] ^ x[67];
  assign t[222] = t[263] ^ x[71];
  assign t[223] = t[264] ^ x[73];
  assign t[224] = t[265] ^ x[75];
  assign t[225] = t[266] ^ x[77];
  assign t[226] = t[267] ^ x[79];
  assign t[227] = t[268] ^ x[83];
  assign t[228] = t[269] ^ x[85];
  assign t[229] = t[270] ^ x[88];
  assign t[22] = ~(t[25] ^ t[34]);
  assign t[230] = t[271] ^ x[92];
  assign t[231] = t[272] ^ x[94];
  assign t[232] = t[273] ^ x[96];
  assign t[233] = t[274] ^ x[98];
  assign t[234] = t[275] ^ x[100];
  assign t[235] = t[276] ^ x[102];
  assign t[236] = t[277] ^ x[104];
  assign t[237] = t[278] ^ x[106];
  assign t[238] = t[279] ^ x[108];
  assign t[239] = t[280] ^ x[110];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[240] = t[281] ^ x[112];
  assign t[241] = (x[0] & x[1]);
  assign t[242] = (x[8] & x[9]);
  assign t[243] = (x[11] & x[12]);
  assign t[244] = (x[14] & x[15]);
  assign t[245] = (x[17] & x[18]);
  assign t[246] = (x[20] & x[21]);
  assign t[247] = (x[23] & x[24]);
  assign t[248] = (x[20] & x[26]);
  assign t[249] = (x[20] & x[28]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[32] & x[33]);
  assign t[251] = (x[35] & x[36]);
  assign t[252] = (x[23] & x[38]);
  assign t[253] = (x[23] & x[40]);
  assign t[254] = (x[42] & x[43]);
  assign t[255] = (x[47] & x[48]);
  assign t[256] = (x[50] & x[51]);
  assign t[257] = (x[20] & x[53]);
  assign t[258] = (x[32] & x[55]);
  assign t[259] = (x[32] & x[57]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[260] = (x[59] & x[60]);
  assign t[261] = (x[35] & x[64]);
  assign t[262] = (x[35] & x[66]);
  assign t[263] = (x[23] & x[70]);
  assign t[264] = (x[42] & x[72]);
  assign t[265] = (x[42] & x[74]);
  assign t[266] = (x[47] & x[76]);
  assign t[267] = (x[47] & x[78]);
  assign t[268] = (x[50] & x[82]);
  assign t[269] = (x[50] & x[84]);
  assign t[26] = ~(t[41] ^ t[42]);
  assign t[270] = (x[86] & x[87]);
  assign t[271] = (x[32] & x[91]);
  assign t[272] = (x[59] & x[93]);
  assign t[273] = (x[59] & x[95]);
  assign t[274] = (x[35] & x[97]);
  assign t[275] = (x[42] & x[99]);
  assign t[276] = (x[47] & x[101]);
  assign t[277] = (x[50] & x[103]);
  assign t[278] = (x[86] & x[105]);
  assign t[279] = (x[86] & x[107]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[280] = (x[59] & x[109]);
  assign t[281] = (x[86] & x[111]);
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[29] = ~(t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[205] | t[54]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[37] = ~(t[61] | t[62]);
  assign t[38] = ~(t[37] ^ t[63]);
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[206] | t[66]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[42] = ~(t[69] ^ t[70]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[44] = ~(t[43] ^ t[73]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[47] = ~(t[203]);
  assign t[48] = ~(t[78] | t[79]);
  assign t[49] = ~(t[78] | t[80]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[204] & t[81];
  assign t[51] = ~(t[82]);
  assign t[52] = ~(t[207]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[83] | t[84]);
  assign t[55] = t[203] ? x[31] : x[30];
  assign t[56] = ~(t[85] & t[86]);
  assign t[57] = ~(t[87] | t[88]);
  assign t[58] = ~(t[209] | t[89]);
  assign t[59] = ~(t[90] | t[91]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[92] ^ t[93]);
  assign t[61] = ~(t[94] | t[95]);
  assign t[62] = ~(t[210] | t[96]);
  assign t[63] = ~(t[97] ^ t[98]);
  assign t[64] = ~(t[211]);
  assign t[65] = ~(t[212]);
  assign t[66] = ~(t[99] | t[100]);
  assign t[67] = ~(t[101] | t[102]);
  assign t[68] = ~(t[213] | t[103]);
  assign t[69] = t[104] ? x[46] : x[45];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[107] | t[108]);
  assign t[72] = ~(t[214] | t[109]);
  assign t[73] = ~(t[110] ^ t[111]);
  assign t[74] = ~(t[112] | t[113]);
  assign t[75] = ~(t[215] | t[114]);
  assign t[76] = ~(t[115] | t[116]);
  assign t[77] = ~(t[117] ^ t[118]);
  assign t[78] = ~(t[119]);
  assign t[79] = t[201] ? t[121] : t[120];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[201] ? t[123] : t[122];
  assign t[81] = ~(t[119] | t[201]);
  assign t[82] = ~(t[124] | t[125]);
  assign t[83] = ~(t[216]);
  assign t[84] = ~(t[207] | t[208]);
  assign t[85] = ~(t[126] | t[127]);
  assign t[86] = ~(t[128] | t[49]);
  assign t[87] = ~(t[217]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[129] | t[130]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = ~(t[219] | t[133]);
  assign t[92] = t[104] ? x[63] : x[62];
  assign t[93] = ~(t[134] & t[106]);
  assign t[94] = ~(t[220]);
  assign t[95] = ~(t[221]);
  assign t[96] = ~(t[135] | t[136]);
  assign t[97] = t[203] ? x[69] : x[68];
  assign t[98] = t[137] | t[138];
  assign t[99] = ~(t[222]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[200];
endmodule

module R1ind142(x, y);
 input [121:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[108] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[31];
  assign t[117] = t[162] ^ x[33];
  assign t[118] = t[163] ^ x[36];
  assign t[119] = t[164] ^ x[39];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[44];
  assign t[121] = t[166] ^ x[48];
  assign t[122] = t[167] ^ x[50];
  assign t[123] = t[168] ^ x[53];
  assign t[124] = t[169] ^ x[56];
  assign t[125] = t[170] ^ x[61];
  assign t[126] = t[171] ^ x[65];
  assign t[127] = t[172] ^ x[67];
  assign t[128] = t[173] ^ x[69];
  assign t[129] = t[174] ^ x[71];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[73];
  assign t[131] = t[176] ^ x[76];
  assign t[132] = t[177] ^ x[78];
  assign t[133] = t[178] ^ x[80];
  assign t[134] = t[179] ^ x[82];
  assign t[135] = t[180] ^ x[84];
  assign t[136] = t[181] ^ x[86];
  assign t[137] = t[182] ^ x[88];
  assign t[138] = t[183] ^ x[90];
  assign t[139] = t[184] ^ x[92];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[94];
  assign t[141] = t[186] ^ x[97];
  assign t[142] = t[187] ^ x[99];
  assign t[143] = t[188] ^ x[101];
  assign t[144] = t[189] ^ x[103];
  assign t[145] = t[190] ^ x[105];
  assign t[146] = t[191] ^ x[107];
  assign t[147] = t[192] ^ x[109];
  assign t[148] = t[193] ^ x[111];
  assign t[149] = t[194] ^ x[113];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[115];
  assign t[151] = t[196] ^ x[117];
  assign t[152] = t[197] ^ x[119];
  assign t[153] = t[198] ^ x[121];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[20] & x[30]);
  assign t[162] = (x[20] & x[32]);
  assign t[163] = (x[34] & x[35]);
  assign t[164] = (x[37] & x[38]);
  assign t[165] = (x[42] & x[43]);
  assign t[166] = (x[25] & x[47]);
  assign t[167] = (x[25] & x[49]);
  assign t[168] = (x[51] & x[52]);
  assign t[169] = (x[54] & x[55]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[59] & x[60]);
  assign t[171] = (x[20] & x[64]);
  assign t[172] = (x[34] & x[66]);
  assign t[173] = (x[34] & x[68]);
  assign t[174] = (x[37] & x[70]);
  assign t[175] = (x[37] & x[72]);
  assign t[176] = (x[74] & x[75]);
  assign t[177] = (x[42] & x[77]);
  assign t[178] = (x[42] & x[79]);
  assign t[179] = (x[25] & x[81]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[51] & x[83]);
  assign t[181] = (x[51] & x[85]);
  assign t[182] = (x[54] & x[87]);
  assign t[183] = (x[54] & x[89]);
  assign t[184] = (x[59] & x[91]);
  assign t[185] = (x[59] & x[93]);
  assign t[186] = (x[95] & x[96]);
  assign t[187] = (x[34] & x[98]);
  assign t[188] = (x[37] & x[100]);
  assign t[189] = (x[74] & x[102]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[74] & x[104]);
  assign t[191] = (x[42] & x[106]);
  assign t[192] = (x[51] & x[108]);
  assign t[193] = (x[54] & x[110]);
  assign t[194] = (x[59] & x[112]);
  assign t[195] = (x[95] & x[114]);
  assign t[196] = (x[95] & x[116]);
  assign t[197] = (x[74] & x[118]);
  assign t[198] = (x[95] & x[120]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] ^ t[43];
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = t[60] | t[115];
  assign t[39] = t[61] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[62] & t[63]);
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[71] | t[45]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[74] | t[118];
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = t[77] | t[119];
  assign t[53] = t[48] ? x[41] : x[40];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[80] & t[81]);
  assign t[56] = t[82] | t[120];
  assign t[57] = t[61] ? x[46] : x[45];
  assign t[58] = ~(t[121]);
  assign t[59] = ~(t[122]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[83] | t[58]);
  assign t[61] = ~(t[24]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[123];
  assign t[64] = ~(t[87] & t[88]);
  assign t[65] = t[89] | t[124];
  assign t[66] = t[61] ? x[58] : x[57];
  assign t[67] = ~(t[90] & t[91]);
  assign t[68] = t[92] | t[125];
  assign t[69] = t[61] ? x[63] : x[62];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[93] & t[94]);
  assign t[71] = ~(t[126]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[128]);
  assign t[74] = ~(t[95] | t[72]);
  assign t[75] = ~(t[129]);
  assign t[76] = ~(t[130]);
  assign t[77] = ~(t[96] | t[75]);
  assign t[78] = ~(t[97] & t[98]);
  assign t[79] = t[99] | t[131];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[132]);
  assign t[81] = ~(t[133]);
  assign t[82] = ~(t[100] | t[80]);
  assign t[83] = ~(t[134]);
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[101] | t[84]);
  assign t[87] = ~(t[137]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[102] | t[87]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[139]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[103] | t[90]);
  assign t[93] = ~(t[104] & t[105]);
  assign t[94] = t[106] | t[141];
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[107] | t[97]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind143(x, y);
 input [121:0] x;
 output y;

 wire [208:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[155]);
  assign t[103] = ~(t[115] & t[116]);
  assign t[104] = ~(t[143] & t[142]);
  assign t[105] = ~(t[156]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[117] & t[118]);
  assign t[115] = ~(t[155] & t[154]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[161] & t[160]);
  assign t[118] = ~(t[163]);
  assign t[119] = t[164] ^ x[2];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[10];
  assign t[121] = t[166] ^ x[13];
  assign t[122] = t[167] ^ x[16];
  assign t[123] = t[168] ^ x[19];
  assign t[124] = t[169] ^ x[22];
  assign t[125] = t[170] ^ x[27];
  assign t[126] = t[171] ^ x[31];
  assign t[127] = t[172] ^ x[33];
  assign t[128] = t[173] ^ x[36];
  assign t[129] = t[174] ^ x[39];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[44];
  assign t[131] = t[176] ^ x[48];
  assign t[132] = t[177] ^ x[50];
  assign t[133] = t[178] ^ x[53];
  assign t[134] = t[179] ^ x[56];
  assign t[135] = t[180] ^ x[61];
  assign t[136] = t[181] ^ x[65];
  assign t[137] = t[182] ^ x[67];
  assign t[138] = t[183] ^ x[69];
  assign t[139] = t[184] ^ x[71];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[73];
  assign t[141] = t[186] ^ x[76];
  assign t[142] = t[187] ^ x[78];
  assign t[143] = t[188] ^ x[80];
  assign t[144] = t[189] ^ x[82];
  assign t[145] = t[190] ^ x[84];
  assign t[146] = t[191] ^ x[86];
  assign t[147] = t[192] ^ x[88];
  assign t[148] = t[193] ^ x[90];
  assign t[149] = t[194] ^ x[92];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[94];
  assign t[151] = t[196] ^ x[97];
  assign t[152] = t[197] ^ x[99];
  assign t[153] = t[198] ^ x[101];
  assign t[154] = t[199] ^ x[103];
  assign t[155] = t[200] ^ x[105];
  assign t[156] = t[201] ^ x[107];
  assign t[157] = t[202] ^ x[109];
  assign t[158] = t[203] ^ x[111];
  assign t[159] = t[204] ^ x[113];
  assign t[15] = ~(t[120] & t[121]);
  assign t[160] = t[205] ^ x[115];
  assign t[161] = t[206] ^ x[117];
  assign t[162] = t[207] ^ x[119];
  assign t[163] = t[208] ^ x[121];
  assign t[164] = (x[0] & x[1]);
  assign t[165] = (x[8] & x[9]);
  assign t[166] = (x[11] & x[12]);
  assign t[167] = (x[14] & x[15]);
  assign t[168] = (x[17] & x[18]);
  assign t[169] = (x[20] & x[21]);
  assign t[16] = ~(t[122] & t[123]);
  assign t[170] = (x[25] & x[26]);
  assign t[171] = (x[20] & x[30]);
  assign t[172] = (x[20] & x[32]);
  assign t[173] = (x[34] & x[35]);
  assign t[174] = (x[37] & x[38]);
  assign t[175] = (x[42] & x[43]);
  assign t[176] = (x[25] & x[47]);
  assign t[177] = (x[25] & x[49]);
  assign t[178] = (x[51] & x[52]);
  assign t[179] = (x[54] & x[55]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[59] & x[60]);
  assign t[181] = (x[20] & x[64]);
  assign t[182] = (x[34] & x[66]);
  assign t[183] = (x[34] & x[68]);
  assign t[184] = (x[37] & x[70]);
  assign t[185] = (x[37] & x[72]);
  assign t[186] = (x[74] & x[75]);
  assign t[187] = (x[42] & x[77]);
  assign t[188] = (x[42] & x[79]);
  assign t[189] = (x[25] & x[81]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[51] & x[83]);
  assign t[191] = (x[51] & x[85]);
  assign t[192] = (x[54] & x[87]);
  assign t[193] = (x[54] & x[89]);
  assign t[194] = (x[59] & x[91]);
  assign t[195] = (x[59] & x[93]);
  assign t[196] = (x[95] & x[96]);
  assign t[197] = (x[34] & x[98]);
  assign t[198] = (x[37] & x[100]);
  assign t[199] = (x[74] & x[102]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[74] & x[104]);
  assign t[201] = (x[42] & x[106]);
  assign t[202] = (x[51] & x[108]);
  assign t[203] = (x[54] & x[110]);
  assign t[204] = (x[59] & x[112]);
  assign t[205] = (x[95] & x[114]);
  assign t[206] = (x[95] & x[116]);
  assign t[207] = (x[74] & x[118]);
  assign t[208] = (x[95] & x[120]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[122]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] & t[124]);
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] ^ t[43];
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = ~(t[60] & t[125]);
  assign t[39] = t[61] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[62] & t[63]);
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = t[69] ^ t[70];
  assign t[45] = ~(t[126]);
  assign t[46] = ~(t[127]);
  assign t[47] = ~(t[71] & t[72]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[75] & t[128]);
  assign t[51] = ~(t[76] & t[77]);
  assign t[52] = ~(t[78] & t[129]);
  assign t[53] = t[48] ? x[41] : x[40];
  assign t[54] = ~(t[79] & t[80]);
  assign t[55] = ~(t[81] & t[82]);
  assign t[56] = ~(t[83] & t[130]);
  assign t[57] = t[17] ? x[46] : x[45];
  assign t[58] = ~(t[131]);
  assign t[59] = ~(t[132]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = ~(t[24]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[133]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[134]);
  assign t[66] = t[61] ? x[58] : x[57];
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = ~(t[94] & t[135]);
  assign t[69] = t[61] ? x[63] : x[62];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[95] & t[96]);
  assign t[71] = ~(t[127] & t[126]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[97] & t[98]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[101] & t[102]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[103] & t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[104] & t[105]);
  assign t[84] = ~(t[132] & t[131]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[147]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[108] & t[109]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[150]);
  assign t[94] = ~(t[110] & t[111]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[114] & t[151]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[119];
endmodule

module R1ind144(x, y);
 input [101:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[135] ^ x[10];
  assign t[101] = t[136] ^ x[13];
  assign t[102] = t[137] ^ x[16];
  assign t[103] = t[138] ^ x[19];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[24];
  assign t[106] = t[141] ^ x[29];
  assign t[107] = t[142] ^ x[31];
  assign t[108] = t[143] ^ x[35];
  assign t[109] = t[144] ^ x[38];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] ^ x[40];
  assign t[111] = t[146] ^ x[43];
  assign t[112] = t[147] ^ x[45];
  assign t[113] = t[148] ^ x[50];
  assign t[114] = t[149] ^ x[52];
  assign t[115] = t[150] ^ x[56];
  assign t[116] = t[151] ^ x[59];
  assign t[117] = t[152] ^ x[61];
  assign t[118] = t[153] ^ x[64];
  assign t[119] = t[154] ^ x[66];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[155] ^ x[71];
  assign t[121] = t[156] ^ x[73];
  assign t[122] = t[157] ^ x[77];
  assign t[123] = t[158] ^ x[79];
  assign t[124] = t[159] ^ x[82];
  assign t[125] = t[160] ^ x[84];
  assign t[126] = t[161] ^ x[86];
  assign t[127] = t[162] ^ x[88];
  assign t[128] = t[163] ^ x[90];
  assign t[129] = t[164] ^ x[93];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[165] ^ x[95];
  assign t[131] = t[166] ^ x[97];
  assign t[132] = t[167] ^ x[99];
  assign t[133] = t[168] ^ x[101];
  assign t[134] = (x[0] & x[1]);
  assign t[135] = (x[8] & x[9]);
  assign t[136] = (x[11] & x[12]);
  assign t[137] = (x[14] & x[15]);
  assign t[138] = (x[17] & x[18]);
  assign t[139] = (x[20] & x[21]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[20] & x[23]);
  assign t[141] = (x[27] & x[28]);
  assign t[142] = (x[27] & x[30]);
  assign t[143] = (x[20] & x[34]);
  assign t[144] = (x[36] & x[37]);
  assign t[145] = (x[36] & x[39]);
  assign t[146] = (x[41] & x[42]);
  assign t[147] = (x[41] & x[44]);
  assign t[148] = (x[48] & x[49]);
  assign t[149] = (x[48] & x[51]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[27] & x[55]);
  assign t[151] = (x[57] & x[58]);
  assign t[152] = (x[57] & x[60]);
  assign t[153] = (x[62] & x[63]);
  assign t[154] = (x[62] & x[65]);
  assign t[155] = (x[69] & x[70]);
  assign t[156] = (x[69] & x[72]);
  assign t[157] = (x[36] & x[76]);
  assign t[158] = (x[41] & x[78]);
  assign t[159] = (x[80] & x[81]);
  assign t[15] = ~(t[100] & t[101]);
  assign t[160] = (x[80] & x[83]);
  assign t[161] = (x[48] & x[85]);
  assign t[162] = (x[57] & x[87]);
  assign t[163] = (x[62] & x[89]);
  assign t[164] = (x[91] & x[92]);
  assign t[165] = (x[91] & x[94]);
  assign t[166] = (x[69] & x[96]);
  assign t[167] = (x[80] & x[98]);
  assign t[168] = (x[91] & x[100]);
  assign t[16] = ~(t[102] & t[103]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = t[47] ? x[26] : x[25];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = t[56] ^ t[41];
  assign t[37] = ~(t[106] & t[57]);
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = t[59] ? x[33] : x[32];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[43];
  assign t[45] = ~(t[108]);
  assign t[46] = ~(t[108] & t[69]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[109] & t[70]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = t[59] ? x[47] : x[46];
  assign t[53] = ~(t[74] & t[75]);
  assign t[54] = ~(t[113] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = t[47] ? x[54] : x[53];
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[24]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[116] & t[79]);
  assign t[61] = ~(t[117] & t[80]);
  assign t[62] = ~(t[118] & t[81]);
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = t[59] ? x[68] : x[67];
  assign t[65] = ~(t[83] & t[84]);
  assign t[66] = ~(t[120] & t[85]);
  assign t[67] = ~(t[121] & t[86]);
  assign t[68] = t[59] ? x[75] : x[74];
  assign t[69] = ~(t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[123]);
  assign t[73] = ~(t[123] & t[88]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126]);
  assign t[77] = ~(t[126] & t[91]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[127]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[127] & t[92]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130] & t[95]);
  assign t[85] = ~(t[131]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[132] & t[97]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[118]);
  assign t[94] = ~(t[133]);
  assign t[95] = ~(t[133] & t[98]);
  assign t[96] = ~(t[120]);
  assign t[97] = ~(t[124]);
  assign t[98] = ~(t[129]);
  assign t[99] = t[134] ^ x[2];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind145(x, y);
 input [121:0] x;
 output y;

 wire [299:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[143] | t[144]);
  assign t[101] = ~(t[145] | t[146]);
  assign t[102] = ~(t[234] | t[147]);
  assign t[103] = t[90] ? x[76] : x[75];
  assign t[104] = ~(t[148] & t[149]);
  assign t[105] = ~(t[235]);
  assign t[106] = ~(t[222] | t[223]);
  assign t[107] = ~(t[236]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[150] | t[151]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[48]);
  assign t[111] = ~(t[136] | t[152]);
  assign t[112] = ~(t[153] | t[154]);
  assign t[113] = ~(t[238]);
  assign t[114] = ~(t[239]);
  assign t[115] = ~(t[155] | t[156]);
  assign t[116] = t[110] ? x[88] : x[87];
  assign t[117] = ~(t[157] & t[158]);
  assign t[118] = ~(t[240]);
  assign t[119] = ~(t[241]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[159] | t[160]);
  assign t[121] = ~(t[161] | t[162]);
  assign t[122] = ~(t[242] | t[163]);
  assign t[123] = t[110] ? x[97] : x[96];
  assign t[124] = ~(t[83] & t[148]);
  assign t[125] = ~(t[213]);
  assign t[126] = ~(t[164] & t[165]);
  assign t[127] = ~(x[4] & t[166]);
  assign t[128] = ~(t[80] | t[167]);
  assign t[129] = ~(t[141] & t[168]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[125] | t[169]);
  assign t[131] = ~(t[125] | t[170]);
  assign t[132] = ~(t[171] & t[214]);
  assign t[133] = ~(t[172] & t[165]);
  assign t[134] = ~(t[243]);
  assign t[135] = ~(t[228] | t[229]);
  assign t[136] = ~(t[80] | t[173]);
  assign t[137] = t[174] | t[175];
  assign t[138] = ~(t[176] & t[177]);
  assign t[139] = ~(t[244]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[230] | t[231]);
  assign t[141] = ~(t[178] | t[179]);
  assign t[142] = ~(t[180] | t[181]);
  assign t[143] = ~(t[245]);
  assign t[144] = ~(t[232] | t[233]);
  assign t[145] = ~(t[246]);
  assign t[146] = ~(t[247]);
  assign t[147] = ~(t[182] | t[183]);
  assign t[148] = ~(t[129] | t[184]);
  assign t[149] = ~(t[128] | t[152]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[248]);
  assign t[151] = ~(t[236] | t[237]);
  assign t[152] = ~(t[80] | t[185]);
  assign t[153] = t[214] & t[186];
  assign t[154] = ~(t[83]);
  assign t[155] = ~(t[249]);
  assign t[156] = ~(t[238] | t[239]);
  assign t[157] = ~(t[178] | t[131]);
  assign t[158] = ~(t[187] | t[175]);
  assign t[159] = ~(t[250]);
  assign t[15] = ~(t[211] & t[212]);
  assign t[160] = ~(t[240] | t[241]);
  assign t[161] = ~(t[251]);
  assign t[162] = ~(t[252]);
  assign t[163] = ~(t[188] | t[189]);
  assign t[164] = ~(x[4] | t[190]);
  assign t[165] = ~(t[214]);
  assign t[166] = ~(t[212] | t[165]);
  assign t[167] = t[211] ? t[132] : t[133];
  assign t[168] = ~(t[125] & t[191]);
  assign t[169] = t[211] ? t[192] : t[133];
  assign t[16] = ~(t[213] & t[214]);
  assign t[170] = t[211] ? t[126] : t[193];
  assign t[171] = x[4] & t[212];
  assign t[172] = ~(x[4] | t[212]);
  assign t[173] = t[211] ? t[193] : t[194];
  assign t[174] = ~(t[83] & t[195]);
  assign t[175] = ~(t[80] | t[196]);
  assign t[176] = ~(t[197] | t[49]);
  assign t[177] = t[125] | t[198];
  assign t[178] = ~(t[125] | t[199]);
  assign t[179] = ~(t[80] | t[200]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[80] | t[201]);
  assign t[181] = ~(t[149] & t[177]);
  assign t[182] = ~(t[253]);
  assign t[183] = ~(t[246] | t[247]);
  assign t[184] = ~(t[202] & t[177]);
  assign t[185] = t[211] ? t[192] : t[203];
  assign t[186] = ~(t[125] | t[211]);
  assign t[187] = ~(t[204]);
  assign t[188] = ~(t[254]);
  assign t[189] = ~(t[251] | t[252]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[212]);
  assign t[191] = ~(t[193] & t[194]);
  assign t[192] = ~(t[171] & t[165]);
  assign t[193] = ~(x[4] & t[205]);
  assign t[194] = ~(t[214] & t[164]);
  assign t[195] = ~(t[166] & t[206]);
  assign t[196] = t[211] ? t[194] : t[193];
  assign t[197] = ~(t[207]);
  assign t[198] = t[211] ? t[193] : t[126];
  assign t[199] = t[211] ? t[133] : t[192];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[211] ? t[126] : t[127];
  assign t[201] = t[211] ? t[203] : t[192];
  assign t[202] = ~(t[153] & t[208]);
  assign t[203] = ~(t[172] & t[214]);
  assign t[204] = ~(t[49] | t[152]);
  assign t[205] = ~(t[212] | t[214]);
  assign t[206] = t[80] & t[211];
  assign t[207] = ~(t[186] & t[209]);
  assign t[208] = t[172] | t[171];
  assign t[209] = ~(t[194] & t[127]);
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[255] ^ x[2];
  assign t[211] = t[256] ^ x[10];
  assign t[212] = t[257] ^ x[13];
  assign t[213] = t[258] ^ x[16];
  assign t[214] = t[259] ^ x[19];
  assign t[215] = t[260] ^ x[22];
  assign t[216] = t[261] ^ x[25];
  assign t[217] = t[262] ^ x[27];
  assign t[218] = t[263] ^ x[29];
  assign t[219] = t[264] ^ x[32];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[37];
  assign t[221] = t[266] ^ x[40];
  assign t[222] = t[267] ^ x[42];
  assign t[223] = t[268] ^ x[44];
  assign t[224] = t[269] ^ x[47];
  assign t[225] = t[270] ^ x[52];
  assign t[226] = t[271] ^ x[55];
  assign t[227] = t[272] ^ x[57];
  assign t[228] = t[273] ^ x[59];
  assign t[229] = t[274] ^ x[61];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[63];
  assign t[231] = t[276] ^ x[65];
  assign t[232] = t[277] ^ x[69];
  assign t[233] = t[278] ^ x[71];
  assign t[234] = t[279] ^ x[74];
  assign t[235] = t[280] ^ x[78];
  assign t[236] = t[281] ^ x[80];
  assign t[237] = t[282] ^ x[82];
  assign t[238] = t[283] ^ x[84];
  assign t[239] = t[284] ^ x[86];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[90];
  assign t[241] = t[286] ^ x[92];
  assign t[242] = t[287] ^ x[95];
  assign t[243] = t[288] ^ x[99];
  assign t[244] = t[289] ^ x[101];
  assign t[245] = t[290] ^ x[103];
  assign t[246] = t[291] ^ x[105];
  assign t[247] = t[292] ^ x[107];
  assign t[248] = t[293] ^ x[109];
  assign t[249] = t[294] ^ x[111];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = t[295] ^ x[113];
  assign t[251] = t[296] ^ x[115];
  assign t[252] = t[297] ^ x[117];
  assign t[253] = t[298] ^ x[119];
  assign t[254] = t[299] ^ x[121];
  assign t[255] = (x[0] & x[1]);
  assign t[256] = (x[8] & x[9]);
  assign t[257] = (x[11] & x[12]);
  assign t[258] = (x[14] & x[15]);
  assign t[259] = (x[17] & x[18]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[20] & x[21]);
  assign t[261] = (x[23] & x[24]);
  assign t[262] = (x[20] & x[26]);
  assign t[263] = (x[20] & x[28]);
  assign t[264] = (x[30] & x[31]);
  assign t[265] = (x[35] & x[36]);
  assign t[266] = (x[38] & x[39]);
  assign t[267] = (x[23] & x[41]);
  assign t[268] = (x[23] & x[43]);
  assign t[269] = (x[45] & x[46]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[50] & x[51]);
  assign t[271] = (x[53] & x[54]);
  assign t[272] = (x[20] & x[56]);
  assign t[273] = (x[30] & x[58]);
  assign t[274] = (x[30] & x[60]);
  assign t[275] = (x[35] & x[62]);
  assign t[276] = (x[35] & x[64]);
  assign t[277] = (x[38] & x[68]);
  assign t[278] = (x[38] & x[70]);
  assign t[279] = (x[72] & x[73]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[23] & x[77]);
  assign t[281] = (x[45] & x[79]);
  assign t[282] = (x[45] & x[81]);
  assign t[283] = (x[50] & x[83]);
  assign t[284] = (x[50] & x[85]);
  assign t[285] = (x[53] & x[89]);
  assign t[286] = (x[53] & x[91]);
  assign t[287] = (x[93] & x[94]);
  assign t[288] = (x[30] & x[98]);
  assign t[289] = (x[35] & x[100]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[290] = (x[38] & x[102]);
  assign t[291] = (x[72] & x[104]);
  assign t[292] = (x[72] & x[106]);
  assign t[293] = (x[45] & x[108]);
  assign t[294] = (x[50] & x[110]);
  assign t[295] = (x[53] & x[112]);
  assign t[296] = (x[93] & x[114]);
  assign t[297] = (x[93] & x[116]);
  assign t[298] = (x[72] & x[118]);
  assign t[299] = (x[93] & x[120]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[215] | t[54]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[36] = ~(t[59] | t[60]);
  assign t[37] = ~(t[46] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[64] ^ t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[66] | t[67]);
  assign t[41] = ~(t[216] | t[68]);
  assign t[42] = ~(t[69] | t[70]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[45] = ~(t[44] ^ t[75]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[47] = ~(t[78] ^ t[79]);
  assign t[48] = ~(t[213]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[82] & t[83]);
  assign t[51] = ~(t[80] | t[84]);
  assign t[52] = ~(t[217]);
  assign t[53] = ~(t[218]);
  assign t[54] = ~(t[85] | t[86]);
  assign t[55] = ~(t[87] | t[88]);
  assign t[56] = ~(t[219] | t[89]);
  assign t[57] = t[90] ? x[34] : x[33];
  assign t[58] = ~(t[91] & t[92]);
  assign t[59] = ~(t[93] | t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[220] | t[95]);
  assign t[61] = ~(t[96] ^ t[97]);
  assign t[62] = ~(t[98] | t[99]);
  assign t[63] = ~(t[221] | t[100]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[65] = ~(t[103] ^ t[104]);
  assign t[66] = ~(t[222]);
  assign t[67] = ~(t[223]);
  assign t[68] = ~(t[105] | t[106]);
  assign t[69] = ~(t[107] | t[108]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[224] | t[109]);
  assign t[71] = t[110] ? x[49] : x[48];
  assign t[72] = ~(t[111] & t[112]);
  assign t[73] = ~(t[113] | t[114]);
  assign t[74] = ~(t[225] | t[115]);
  assign t[75] = ~(t[116] ^ t[117]);
  assign t[76] = ~(t[118] | t[119]);
  assign t[77] = ~(t[226] | t[120]);
  assign t[78] = ~(t[121] | t[122]);
  assign t[79] = ~(t[123] ^ t[124]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[125]);
  assign t[81] = t[211] ? t[127] : t[126];
  assign t[82] = ~(t[128] | t[129]);
  assign t[83] = ~(t[130] | t[131]);
  assign t[84] = t[211] ? t[133] : t[132];
  assign t[85] = ~(t[227]);
  assign t[86] = ~(t[217] | t[218]);
  assign t[87] = ~(t[228]);
  assign t[88] = ~(t[229]);
  assign t[89] = ~(t[134] | t[135]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[48]);
  assign t[91] = ~(t[128] | t[136]);
  assign t[92] = ~(t[137] | t[138]);
  assign t[93] = ~(t[230]);
  assign t[94] = ~(t[231]);
  assign t[95] = ~(t[139] | t[140]);
  assign t[96] = t[90] ? x[67] : x[66];
  assign t[97] = ~(t[141] & t[142]);
  assign t[98] = ~(t[232]);
  assign t[99] = ~(t[233]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[210];
endmodule

module R1ind146(x, y);
 input [85:0] x;
 output y;

 wire [142:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[65];
  assign t[101] = t[133] ^ x[67];
  assign t[102] = t[134] ^ x[69];
  assign t[103] = t[135] ^ x[71];
  assign t[104] = t[136] ^ x[73];
  assign t[105] = t[137] ^ x[75];
  assign t[106] = t[138] ^ x[77];
  assign t[107] = t[139] ^ x[79];
  assign t[108] = t[140] ^ x[81];
  assign t[109] = t[141] ^ x[83];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[85];
  assign t[111] = (x[0] & x[1]);
  assign t[112] = (x[8] & x[9]);
  assign t[113] = (x[11] & x[12]);
  assign t[114] = (x[14] & x[15]);
  assign t[115] = (x[17] & x[18]);
  assign t[116] = (x[20] & x[21]);
  assign t[117] = (x[0] & x[23]);
  assign t[118] = (x[20] & x[27]);
  assign t[119] = (x[20] & x[29]);
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = (x[31] & x[32]);
  assign t[121] = (x[36] & x[37]);
  assign t[122] = (x[0] & x[41]);
  assign t[123] = (x[43] & x[44]);
  assign t[124] = (x[20] & x[46]);
  assign t[125] = (x[31] & x[48]);
  assign t[126] = (x[31] & x[50]);
  assign t[127] = (x[52] & x[53]);
  assign t[128] = (x[36] & x[55]);
  assign t[129] = (x[36] & x[57]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[130] = (x[59] & x[60]);
  assign t[131] = (x[0] & x[62]);
  assign t[132] = (x[43] & x[64]);
  assign t[133] = (x[43] & x[66]);
  assign t[134] = (x[31] & x[68]);
  assign t[135] = (x[52] & x[70]);
  assign t[136] = (x[52] & x[72]);
  assign t[137] = (x[36] & x[74]);
  assign t[138] = (x[59] & x[76]);
  assign t[139] = (x[59] & x[78]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = (x[43] & x[80]);
  assign t[141] = (x[52] & x[82]);
  assign t[142] = (x[59] & x[84]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[80] & t[81]);
  assign t[16] = ~(t[82] & t[83]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[82]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[36] & t[37]);
  assign t[27] = t[38] | t[84];
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[43] & t[44]);
  assign t[31] = t[45] ^ t[46];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] | t[85];
  assign t[34] = t[17] ? x[26] : x[25];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = ~(t[86]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[52] | t[36]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[55] | t[88];
  assign t[41] = t[56] ? x[35] : x[34];
  assign t[42] = ~(t[57] & t[58]);
  assign t[43] = ~(t[59] & t[60]);
  assign t[44] = t[61] | t[89];
  assign t[45] = t[56] ? x[40] : x[39];
  assign t[46] = ~(t[62] & t[63]);
  assign t[47] = ~(t[79]);
  assign t[48] = ~(t[90]);
  assign t[49] = ~(t[64] | t[47]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[65] & t[66]);
  assign t[51] = t[67] | t[91];
  assign t[52] = ~(t[92]);
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[68] | t[53]);
  assign t[56] = ~(t[23]);
  assign t[57] = ~(t[69] & t[70]);
  assign t[58] = t[71] | t[95];
  assign t[59] = ~(t[96]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[97]);
  assign t[61] = ~(t[72] | t[59]);
  assign t[62] = ~(t[73] & t[74]);
  assign t[63] = t[75] | t[98];
  assign t[64] = ~(t[99]);
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[76] | t[65]);
  assign t[68] = ~(t[102]);
  assign t[69] = ~(t[103]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[77] | t[69]);
  assign t[72] = ~(t[105]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[78] | t[73]);
  assign t[76] = ~(t[108]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = t[111] ^ x[2];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[112] ^ x[10];
  assign t[81] = t[113] ^ x[13];
  assign t[82] = t[114] ^ x[16];
  assign t[83] = t[115] ^ x[19];
  assign t[84] = t[116] ^ x[22];
  assign t[85] = t[117] ^ x[24];
  assign t[86] = t[118] ^ x[28];
  assign t[87] = t[119] ^ x[30];
  assign t[88] = t[120] ^ x[33];
  assign t[89] = t[121] ^ x[38];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[122] ^ x[42];
  assign t[91] = t[123] ^ x[45];
  assign t[92] = t[124] ^ x[47];
  assign t[93] = t[125] ^ x[49];
  assign t[94] = t[126] ^ x[51];
  assign t[95] = t[127] ^ x[54];
  assign t[96] = t[128] ^ x[56];
  assign t[97] = t[129] ^ x[58];
  assign t[98] = t[130] ^ x[61];
  assign t[99] = t[131] ^ x[63];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[79];
endmodule

module R1ind147(x, y);
 input [85:0] x;
 output y;

 wire [149:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[49];
  assign t[101] = t[133] ^ x[51];
  assign t[102] = t[134] ^ x[53];
  assign t[103] = t[135] ^ x[56];
  assign t[104] = t[136] ^ x[58];
  assign t[105] = t[137] ^ x[60];
  assign t[106] = t[138] ^ x[63];
  assign t[107] = t[139] ^ x[65];
  assign t[108] = t[140] ^ x[67];
  assign t[109] = t[141] ^ x[69];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[71];
  assign t[111] = t[143] ^ x[73];
  assign t[112] = t[144] ^ x[75];
  assign t[113] = t[145] ^ x[77];
  assign t[114] = t[146] ^ x[79];
  assign t[115] = t[147] ^ x[81];
  assign t[116] = t[148] ^ x[83];
  assign t[117] = t[149] ^ x[85];
  assign t[118] = (x[0] & x[1]);
  assign t[119] = (x[8] & x[9]);
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = (x[11] & x[12]);
  assign t[121] = (x[14] & x[15]);
  assign t[122] = (x[17] & x[18]);
  assign t[123] = (x[20] & x[21]);
  assign t[124] = (x[0] & x[23]);
  assign t[125] = (x[20] & x[27]);
  assign t[126] = (x[20] & x[29]);
  assign t[127] = (x[31] & x[32]);
  assign t[128] = (x[36] & x[37]);
  assign t[129] = (x[0] & x[41]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[130] = (x[0] & x[43]);
  assign t[131] = (x[45] & x[46]);
  assign t[132] = (x[20] & x[48]);
  assign t[133] = (x[31] & x[50]);
  assign t[134] = (x[31] & x[52]);
  assign t[135] = (x[54] & x[55]);
  assign t[136] = (x[36] & x[57]);
  assign t[137] = (x[36] & x[59]);
  assign t[138] = (x[61] & x[62]);
  assign t[139] = (x[45] & x[64]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = (x[45] & x[66]);
  assign t[141] = (x[31] & x[68]);
  assign t[142] = (x[54] & x[70]);
  assign t[143] = (x[54] & x[72]);
  assign t[144] = (x[36] & x[74]);
  assign t[145] = (x[61] & x[76]);
  assign t[146] = (x[61] & x[78]);
  assign t[147] = (x[45] & x[80]);
  assign t[148] = (x[54] & x[82]);
  assign t[149] = (x[61] & x[84]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[87] & t[88]);
  assign t[16] = ~(t[89] & t[90]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[89]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[36] & t[37]);
  assign t[27] = ~(t[38] & t[91]);
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[43] & t[44]);
  assign t[31] = t[45] ^ t[46];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = ~(t[49] & t[92]);
  assign t[34] = t[17] ? x[26] : x[25];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = ~(t[93]);
  assign t[37] = ~(t[94]);
  assign t[38] = ~(t[52] & t[53]);
  assign t[39] = ~(t[54] & t[55]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[56] & t[95]);
  assign t[41] = t[57] ? x[35] : x[34];
  assign t[42] = ~(t[58] & t[59]);
  assign t[43] = ~(t[60] & t[61]);
  assign t[44] = ~(t[62] & t[96]);
  assign t[45] = t[57] ? x[40] : x[39];
  assign t[46] = ~(t[63] & t[64]);
  assign t[47] = ~(t[97]);
  assign t[48] = ~(t[98]);
  assign t[49] = ~(t[65] & t[66]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[67] & t[68]);
  assign t[51] = ~(t[69] & t[99]);
  assign t[52] = ~(t[94] & t[93]);
  assign t[53] = ~(t[100]);
  assign t[54] = ~(t[101]);
  assign t[55] = ~(t[102]);
  assign t[56] = ~(t[70] & t[71]);
  assign t[57] = ~(t[23]);
  assign t[58] = ~(t[72] & t[73]);
  assign t[59] = ~(t[74] & t[103]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[104]);
  assign t[61] = ~(t[105]);
  assign t[62] = ~(t[75] & t[76]);
  assign t[63] = ~(t[77] & t[78]);
  assign t[64] = ~(t[79] & t[106]);
  assign t[65] = ~(t[98] & t[97]);
  assign t[66] = ~(t[86]);
  assign t[67] = ~(t[107]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[80] & t[81]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[102] & t[101]);
  assign t[71] = ~(t[109]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[82] & t[83]);
  assign t[75] = ~(t[105] & t[104]);
  assign t[76] = ~(t[112]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[84] & t[85]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[108] & t[107]);
  assign t[81] = ~(t[115]);
  assign t[82] = ~(t[111] & t[110]);
  assign t[83] = ~(t[116]);
  assign t[84] = ~(t[114] & t[113]);
  assign t[85] = ~(t[117]);
  assign t[86] = t[118] ^ x[2];
  assign t[87] = t[119] ^ x[10];
  assign t[88] = t[120] ^ x[13];
  assign t[89] = t[121] ^ x[16];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[122] ^ x[19];
  assign t[91] = t[123] ^ x[22];
  assign t[92] = t[124] ^ x[24];
  assign t[93] = t[125] ^ x[28];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[33];
  assign t[96] = t[128] ^ x[38];
  assign t[97] = t[129] ^ x[42];
  assign t[98] = t[130] ^ x[44];
  assign t[99] = t[131] ^ x[47];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[86];
endmodule

module R1ind148(x, y);
 input [73:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = (x[11] & x[12]);
  assign t[101] = (x[14] & x[15]);
  assign t[102] = (x[17] & x[18]);
  assign t[103] = (x[20] & x[21]);
  assign t[104] = (x[20] & x[23]);
  assign t[105] = (x[0] & x[25]);
  assign t[106] = (x[0] & x[27]);
  assign t[107] = (x[20] & x[31]);
  assign t[108] = (x[33] & x[34]);
  assign t[109] = (x[33] & x[36]);
  assign t[10] = ~(x[3]);
  assign t[110] = (x[40] & x[41]);
  assign t[111] = (x[40] & x[43]);
  assign t[112] = (x[0] & x[47]);
  assign t[113] = (x[49] & x[50]);
  assign t[114] = (x[49] & x[52]);
  assign t[115] = (x[33] & x[54]);
  assign t[116] = (x[56] & x[57]);
  assign t[117] = (x[56] & x[59]);
  assign t[118] = (x[40] & x[61]);
  assign t[119] = (x[63] & x[64]);
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = (x[63] & x[66]);
  assign t[121] = (x[49] & x[68]);
  assign t[122] = (x[56] & x[70]);
  assign t[123] = (x[63] & x[72]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[73] & t[74]);
  assign t[16] = ~(t[75] & t[76]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[75]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[77] & t[36]);
  assign t[27] = ~(t[78] & t[37]);
  assign t[28] = ~(t[38] & t[39]);
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[42] & t[43]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[79] & t[46]);
  assign t[33] = ~(t[80] & t[47]);
  assign t[34] = t[17] ? x[30] : x[29];
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = ~(t[81]);
  assign t[37] = ~(t[81] & t[50]);
  assign t[38] = ~(t[82] & t[51]);
  assign t[39] = ~(t[83] & t[52]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[53] ? x[39] : x[38];
  assign t[41] = ~(t[54] & t[55]);
  assign t[42] = ~(t[84] & t[56]);
  assign t[43] = ~(t[85] & t[57]);
  assign t[44] = t[53] ? x[46] : x[45];
  assign t[45] = ~(t[58] & t[59]);
  assign t[46] = ~(t[86]);
  assign t[47] = ~(t[86] & t[60]);
  assign t[48] = ~(t[87] & t[61]);
  assign t[49] = ~(t[88] & t[62]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[77]);
  assign t[51] = ~(t[89]);
  assign t[52] = ~(t[89] & t[63]);
  assign t[53] = ~(t[23]);
  assign t[54] = ~(t[90] & t[64]);
  assign t[55] = ~(t[91] & t[65]);
  assign t[56] = ~(t[92]);
  assign t[57] = ~(t[92] & t[66]);
  assign t[58] = ~(t[93] & t[67]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[79]);
  assign t[61] = ~(t[95]);
  assign t[62] = ~(t[95] & t[69]);
  assign t[63] = ~(t[82]);
  assign t[64] = ~(t[96]);
  assign t[65] = ~(t[96] & t[70]);
  assign t[66] = ~(t[84]);
  assign t[67] = ~(t[97]);
  assign t[68] = ~(t[97] & t[71]);
  assign t[69] = ~(t[87]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[90]);
  assign t[71] = ~(t[93]);
  assign t[72] = t[98] ^ x[2];
  assign t[73] = t[99] ^ x[10];
  assign t[74] = t[100] ^ x[13];
  assign t[75] = t[101] ^ x[16];
  assign t[76] = t[102] ^ x[19];
  assign t[77] = t[103] ^ x[22];
  assign t[78] = t[104] ^ x[24];
  assign t[79] = t[105] ^ x[26];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[106] ^ x[28];
  assign t[81] = t[107] ^ x[32];
  assign t[82] = t[108] ^ x[35];
  assign t[83] = t[109] ^ x[37];
  assign t[84] = t[110] ^ x[42];
  assign t[85] = t[111] ^ x[44];
  assign t[86] = t[112] ^ x[48];
  assign t[87] = t[113] ^ x[51];
  assign t[88] = t[114] ^ x[53];
  assign t[89] = t[115] ^ x[55];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[116] ^ x[58];
  assign t[91] = t[117] ^ x[60];
  assign t[92] = t[118] ^ x[62];
  assign t[93] = t[119] ^ x[65];
  assign t[94] = t[120] ^ x[67];
  assign t[95] = t[121] ^ x[69];
  assign t[96] = t[122] ^ x[71];
  assign t[97] = t[123] ^ x[73];
  assign t[98] = (x[0] & x[1]);
  assign t[99] = (x[8] & x[9]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[72];
endmodule

module R1ind149(x, y);
 input [85:0] x;
 output y;

 wire [214:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[176]);
  assign t[101] = ~(t[119] | t[120]);
  assign t[102] = ~(t[39]);
  assign t[103] = ~(t[121] | t[122]);
  assign t[104] = ~(t[123] & t[124]);
  assign t[105] = ~(t[177]);
  assign t[106] = ~(t[169] | t[170]);
  assign t[107] = ~(t[178]);
  assign t[108] = ~(t[179]);
  assign t[109] = ~(t[125] | t[126]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[113] | t[127]);
  assign t[111] = ~(t[180]);
  assign t[112] = ~(t[172] | t[173]);
  assign t[113] = ~(t[42] | t[128]);
  assign t[114] = ~(t[129]);
  assign t[115] = ~(t[130] & t[94]);
  assign t[116] = ~(t[131] & t[94]);
  assign t[117] = ~(t[96] & t[94]);
  assign t[118] = ~(t[153]);
  assign t[119] = ~(t[181]);
  assign t[11] = ~(t[17] ^ t[14]);
  assign t[120] = ~(t[175] | t[176]);
  assign t[121] = ~(t[132] & t[41]);
  assign t[122] = t[28] | t[133];
  assign t[123] = t[155] & t[134];
  assign t[124] = t[130] | t[131];
  assign t[125] = ~(t[182]);
  assign t[126] = ~(t[178] | t[179]);
  assign t[127] = ~(t[135] & t[136]);
  assign t[128] = t[152] ? t[137] : t[115];
  assign t[129] = ~(t[138] | t[139]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(x[4] | t[153]);
  assign t[131] = x[4] & t[153];
  assign t[132] = ~(t[134] & t[140]);
  assign t[133] = ~(t[42] | t[141]);
  assign t[134] = ~(t[66] | t[152]);
  assign t[135] = ~(t[142] | t[143]);
  assign t[136] = ~(t[66] & t[144]);
  assign t[137] = ~(t[131] & t[155]);
  assign t[138] = ~(t[42] | t[145]);
  assign t[139] = ~(t[42] | t[146]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = ~(t[68] & t[147]);
  assign t[141] = t[152] ? t[148] : t[116];
  assign t[142] = ~(t[66] | t[149]);
  assign t[143] = ~(t[42] | t[150]);
  assign t[144] = ~(t[67] & t[68]);
  assign t[145] = t[152] ? t[147] : t[117];
  assign t[146] = t[152] ? t[116] : t[148];
  assign t[147] = ~(x[4] & t[64]);
  assign t[148] = ~(t[130] & t[155]);
  assign t[149] = t[152] ? t[115] : t[116];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[152] ? t[117] : t[147];
  assign t[151] = t[183] ^ x[2];
  assign t[152] = t[184] ^ x[10];
  assign t[153] = t[185] ^ x[13];
  assign t[154] = t[186] ^ x[16];
  assign t[155] = t[187] ^ x[19];
  assign t[156] = t[188] ^ x[22];
  assign t[157] = t[189] ^ x[24];
  assign t[158] = t[190] ^ x[26];
  assign t[159] = t[191] ^ x[28];
  assign t[15] = ~(t[152] & t[153]);
  assign t[160] = t[192] ^ x[31];
  assign t[161] = t[193] ^ x[34];
  assign t[162] = t[194] ^ x[36];
  assign t[163] = t[195] ^ x[38];
  assign t[164] = t[196] ^ x[41];
  assign t[165] = t[197] ^ x[45];
  assign t[166] = t[198] ^ x[47];
  assign t[167] = t[199] ^ x[49];
  assign t[168] = t[200] ^ x[52];
  assign t[169] = t[201] ^ x[56];
  assign t[16] = ~(t[154] & t[155]);
  assign t[170] = t[202] ^ x[58];
  assign t[171] = t[203] ^ x[61];
  assign t[172] = t[204] ^ x[65];
  assign t[173] = t[205] ^ x[67];
  assign t[174] = t[206] ^ x[69];
  assign t[175] = t[207] ^ x[71];
  assign t[176] = t[208] ^ x[73];
  assign t[177] = t[209] ^ x[75];
  assign t[178] = t[210] ^ x[77];
  assign t[179] = t[211] ^ x[79];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[212] ^ x[81];
  assign t[181] = t[213] ^ x[83];
  assign t[182] = t[214] ^ x[85];
  assign t[183] = (x[0] & x[1]);
  assign t[184] = (x[8] & x[9]);
  assign t[185] = (x[11] & x[12]);
  assign t[186] = (x[14] & x[15]);
  assign t[187] = (x[17] & x[18]);
  assign t[188] = (x[20] & x[21]);
  assign t[189] = (x[0] & x[23]);
  assign t[18] = t[26] ? x[7] : x[6];
  assign t[190] = (x[20] & x[25]);
  assign t[191] = (x[20] & x[27]);
  assign t[192] = (x[29] & x[30]);
  assign t[193] = (x[32] & x[33]);
  assign t[194] = (x[0] & x[35]);
  assign t[195] = (x[0] & x[37]);
  assign t[196] = (x[39] & x[40]);
  assign t[197] = (x[20] & x[44]);
  assign t[198] = (x[29] & x[46]);
  assign t[199] = (x[29] & x[48]);
  assign t[19] = t[27] | t[28];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[50] & x[51]);
  assign t[201] = (x[32] & x[55]);
  assign t[202] = (x[32] & x[57]);
  assign t[203] = (x[59] & x[60]);
  assign t[204] = (x[39] & x[64]);
  assign t[205] = (x[39] & x[66]);
  assign t[206] = (x[29] & x[68]);
  assign t[207] = (x[50] & x[70]);
  assign t[208] = (x[50] & x[72]);
  assign t[209] = (x[32] & x[74]);
  assign t[20] = ~(t[29] | t[30]);
  assign t[210] = (x[59] & x[76]);
  assign t[211] = (x[59] & x[78]);
  assign t[212] = (x[39] & x[80]);
  assign t[213] = (x[50] & x[82]);
  assign t[214] = (x[59] & x[84]);
  assign t[21] = ~(t[24] ^ t[12]);
  assign t[22] = x[4] ? t[32] : t[31];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[24] = ~(t[35] | t[36]);
  assign t[25] = ~(t[37] ^ t[38]);
  assign t[26] = ~(t[39]);
  assign t[27] = ~(t[40] & t[41]);
  assign t[28] = ~(t[42] | t[43]);
  assign t[29] = ~(t[44] | t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[156] | t[46]);
  assign t[31] = ~(t[47] | t[48]);
  assign t[32] = ~(t[49] ^ t[50]);
  assign t[33] = ~(t[51] | t[52]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[157] | t[57]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = ~(t[60] ^ t[61]);
  assign t[39] = ~(t[154]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[62] | t[63]);
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = ~(t[66]);
  assign t[43] = t[152] ? t[68] : t[67];
  assign t[44] = ~(t[158]);
  assign t[45] = ~(t[159]);
  assign t[46] = ~(t[69] | t[70]);
  assign t[47] = ~(t[71] | t[72]);
  assign t[48] = ~(t[160] | t[73]);
  assign t[49] = ~(t[74] | t[75]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[76] ^ t[77]);
  assign t[51] = ~(t[78] | t[79]);
  assign t[52] = ~(t[161] | t[80]);
  assign t[53] = ~(t[81] | t[82]);
  assign t[54] = ~(t[83] ^ t[84]);
  assign t[55] = ~(t[162]);
  assign t[56] = ~(t[163]);
  assign t[57] = ~(t[85] | t[86]);
  assign t[58] = ~(t[87] | t[88]);
  assign t[59] = ~(t[164] | t[89]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[26] ? x[43] : x[42];
  assign t[61] = ~(t[90] & t[91]);
  assign t[62] = ~(t[66] | t[92]);
  assign t[63] = ~(t[66] | t[93]);
  assign t[64] = ~(t[153] | t[94]);
  assign t[65] = t[42] & t[152];
  assign t[66] = ~(t[154]);
  assign t[67] = ~(x[4] & t[95]);
  assign t[68] = ~(t[155] & t[96]);
  assign t[69] = ~(t[165]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[158] | t[159]);
  assign t[71] = ~(t[166]);
  assign t[72] = ~(t[167]);
  assign t[73] = ~(t[97] | t[98]);
  assign t[74] = ~(t[99] | t[100]);
  assign t[75] = ~(t[168] | t[101]);
  assign t[76] = t[102] ? x[54] : x[53];
  assign t[77] = ~(t[103] & t[104]);
  assign t[78] = ~(t[169]);
  assign t[79] = ~(t[170]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[105] | t[106]);
  assign t[81] = ~(t[107] | t[108]);
  assign t[82] = ~(t[171] | t[109]);
  assign t[83] = t[102] ? x[63] : x[62];
  assign t[84] = ~(t[110] & t[41]);
  assign t[85] = ~(t[151]);
  assign t[86] = ~(t[162] | t[163]);
  assign t[87] = ~(t[172]);
  assign t[88] = ~(t[173]);
  assign t[89] = ~(t[111] | t[112]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[113]);
  assign t[91] = ~(t[114] | t[28]);
  assign t[92] = t[152] ? t[116] : t[115];
  assign t[93] = t[152] ? t[117] : t[67];
  assign t[94] = ~(t[155]);
  assign t[95] = ~(t[153] | t[155]);
  assign t[96] = ~(x[4] | t[118]);
  assign t[97] = ~(t[174]);
  assign t[98] = ~(t[166] | t[167]);
  assign t[99] = ~(t[175]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[151];
endmodule

module R1ind150(x, y);
 input [121:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[107] | t[100]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[108] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[31];
  assign t[117] = t[162] ^ x[33];
  assign t[118] = t[163] ^ x[36];
  assign t[119] = t[164] ^ x[39];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[44];
  assign t[121] = t[166] ^ x[48];
  assign t[122] = t[167] ^ x[50];
  assign t[123] = t[168] ^ x[53];
  assign t[124] = t[169] ^ x[56];
  assign t[125] = t[170] ^ x[61];
  assign t[126] = t[171] ^ x[65];
  assign t[127] = t[172] ^ x[67];
  assign t[128] = t[173] ^ x[69];
  assign t[129] = t[174] ^ x[71];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[73];
  assign t[131] = t[176] ^ x[75];
  assign t[132] = t[177] ^ x[77];
  assign t[133] = t[178] ^ x[79];
  assign t[134] = t[179] ^ x[81];
  assign t[135] = t[180] ^ x[83];
  assign t[136] = t[181] ^ x[85];
  assign t[137] = t[182] ^ x[87];
  assign t[138] = t[183] ^ x[90];
  assign t[139] = t[184] ^ x[92];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[94];
  assign t[141] = t[186] ^ x[97];
  assign t[142] = t[187] ^ x[99];
  assign t[143] = t[188] ^ x[101];
  assign t[144] = t[189] ^ x[103];
  assign t[145] = t[190] ^ x[105];
  assign t[146] = t[191] ^ x[107];
  assign t[147] = t[192] ^ x[109];
  assign t[148] = t[193] ^ x[111];
  assign t[149] = t[194] ^ x[113];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[115];
  assign t[151] = t[196] ^ x[117];
  assign t[152] = t[197] ^ x[119];
  assign t[153] = t[198] ^ x[121];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[20] & x[30]);
  assign t[162] = (x[20] & x[32]);
  assign t[163] = (x[34] & x[35]);
  assign t[164] = (x[37] & x[38]);
  assign t[165] = (x[42] & x[43]);
  assign t[166] = (x[25] & x[47]);
  assign t[167] = (x[25] & x[49]);
  assign t[168] = (x[51] & x[52]);
  assign t[169] = (x[54] & x[55]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[59] & x[60]);
  assign t[171] = (x[20] & x[64]);
  assign t[172] = (x[34] & x[66]);
  assign t[173] = (x[34] & x[68]);
  assign t[174] = (x[37] & x[70]);
  assign t[175] = (x[37] & x[72]);
  assign t[176] = (x[42] & x[74]);
  assign t[177] = (x[42] & x[76]);
  assign t[178] = (x[25] & x[78]);
  assign t[179] = (x[51] & x[80]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[51] & x[82]);
  assign t[181] = (x[54] & x[84]);
  assign t[182] = (x[54] & x[86]);
  assign t[183] = (x[88] & x[89]);
  assign t[184] = (x[59] & x[91]);
  assign t[185] = (x[59] & x[93]);
  assign t[186] = (x[95] & x[96]);
  assign t[187] = (x[34] & x[98]);
  assign t[188] = (x[37] & x[100]);
  assign t[189] = (x[42] & x[102]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[51] & x[104]);
  assign t[191] = (x[54] & x[106]);
  assign t[192] = (x[88] & x[108]);
  assign t[193] = (x[88] & x[110]);
  assign t[194] = (x[59] & x[112]);
  assign t[195] = (x[95] & x[114]);
  assign t[196] = (x[95] & x[116]);
  assign t[197] = (x[88] & x[118]);
  assign t[198] = (x[95] & x[120]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[33];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[41];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = t[58] | t[115];
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[68];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[69] | t[45]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = t[72] | t[118];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = t[75] | t[119];
  assign t[52] = t[76] ? x[41] : x[40];
  assign t[53] = ~(t[77] & t[78]);
  assign t[54] = t[79] | t[120];
  assign t[55] = t[76] ? x[46] : x[45];
  assign t[56] = ~(t[121]);
  assign t[57] = ~(t[122]);
  assign t[58] = ~(t[80] | t[56]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[83] | t[123];
  assign t[61] = ~(t[84] & t[85]);
  assign t[62] = t[86] | t[124];
  assign t[63] = t[87] ? x[58] : x[57];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = t[92] | t[125];
  assign t[67] = t[87] ? x[63] : x[62];
  assign t[68] = ~(t[93] & t[94]);
  assign t[69] = ~(t[126]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[128]);
  assign t[72] = ~(t[95] | t[70]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[96] | t[73]);
  assign t[76] = ~(t[24]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[97] | t[77]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[98] | t[81]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[99] | t[84]);
  assign t[87] = ~(t[24]);
  assign t[88] = ~(t[100] & t[101]);
  assign t[89] = t[102] | t[138];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[139]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[103] | t[90]);
  assign t[93] = ~(t[104] & t[105]);
  assign t[94] = t[106] | t[141];
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind151(x, y);
 input [121:0] x;
 output y;

 wire [206:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[152]);
  assign t[101] = ~(t[143] & t[142]);
  assign t[102] = ~(t[153]);
  assign t[103] = ~(t[145] & t[144]);
  assign t[104] = ~(t[154]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[113] & t[114]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[157]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[115] & t[116]);
  assign t[113] = ~(t[156] & t[155]);
  assign t[114] = ~(t[160]);
  assign t[115] = ~(t[159] & t[158]);
  assign t[116] = ~(t[161]);
  assign t[117] = t[162] ^ x[2];
  assign t[118] = t[163] ^ x[8];
  assign t[119] = t[164] ^ x[11];
  assign t[11] = t[15] ? x[19] : x[18];
  assign t[120] = t[165] ^ x[14];
  assign t[121] = t[166] ^ x[17];
  assign t[122] = t[167] ^ x[22];
  assign t[123] = t[168] ^ x[27];
  assign t[124] = t[169] ^ x[31];
  assign t[125] = t[170] ^ x[33];
  assign t[126] = t[171] ^ x[36];
  assign t[127] = t[172] ^ x[39];
  assign t[128] = t[173] ^ x[44];
  assign t[129] = t[174] ^ x[48];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[175] ^ x[50];
  assign t[131] = t[176] ^ x[53];
  assign t[132] = t[177] ^ x[56];
  assign t[133] = t[178] ^ x[61];
  assign t[134] = t[179] ^ x[65];
  assign t[135] = t[180] ^ x[67];
  assign t[136] = t[181] ^ x[69];
  assign t[137] = t[182] ^ x[71];
  assign t[138] = t[183] ^ x[73];
  assign t[139] = t[184] ^ x[75];
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = t[185] ^ x[77];
  assign t[141] = t[186] ^ x[79];
  assign t[142] = t[187] ^ x[81];
  assign t[143] = t[188] ^ x[83];
  assign t[144] = t[189] ^ x[85];
  assign t[145] = t[190] ^ x[87];
  assign t[146] = t[191] ^ x[90];
  assign t[147] = t[192] ^ x[92];
  assign t[148] = t[193] ^ x[94];
  assign t[149] = t[194] ^ x[97];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[195] ^ x[99];
  assign t[151] = t[196] ^ x[101];
  assign t[152] = t[197] ^ x[103];
  assign t[153] = t[198] ^ x[105];
  assign t[154] = t[199] ^ x[107];
  assign t[155] = t[200] ^ x[109];
  assign t[156] = t[201] ^ x[111];
  assign t[157] = t[202] ^ x[113];
  assign t[158] = t[203] ^ x[115];
  assign t[159] = t[204] ^ x[117];
  assign t[15] = ~(t[22]);
  assign t[160] = t[205] ^ x[119];
  assign t[161] = t[206] ^ x[121];
  assign t[162] = (x[0] & x[1]);
  assign t[163] = (x[6] & x[7]);
  assign t[164] = (x[9] & x[10]);
  assign t[165] = (x[12] & x[13]);
  assign t[166] = (x[15] & x[16]);
  assign t[167] = (x[20] & x[21]);
  assign t[168] = (x[25] & x[26]);
  assign t[169] = (x[20] & x[30]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[170] = (x[20] & x[32]);
  assign t[171] = (x[34] & x[35]);
  assign t[172] = (x[37] & x[38]);
  assign t[173] = (x[42] & x[43]);
  assign t[174] = (x[25] & x[47]);
  assign t[175] = (x[25] & x[49]);
  assign t[176] = (x[51] & x[52]);
  assign t[177] = (x[54] & x[55]);
  assign t[178] = (x[59] & x[60]);
  assign t[179] = (x[20] & x[64]);
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[180] = (x[34] & x[66]);
  assign t[181] = (x[34] & x[68]);
  assign t[182] = (x[37] & x[70]);
  assign t[183] = (x[37] & x[72]);
  assign t[184] = (x[42] & x[74]);
  assign t[185] = (x[42] & x[76]);
  assign t[186] = (x[25] & x[78]);
  assign t[187] = (x[51] & x[80]);
  assign t[188] = (x[51] & x[82]);
  assign t[189] = (x[54] & x[84]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[190] = (x[54] & x[86]);
  assign t[191] = (x[88] & x[89]);
  assign t[192] = (x[59] & x[91]);
  assign t[193] = (x[59] & x[93]);
  assign t[194] = (x[95] & x[96]);
  assign t[195] = (x[34] & x[98]);
  assign t[196] = (x[37] & x[100]);
  assign t[197] = (x[42] & x[102]);
  assign t[198] = (x[51] & x[104]);
  assign t[199] = (x[54] & x[106]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[200] = (x[88] & x[108]);
  assign t[201] = (x[88] & x[110]);
  assign t[202] = (x[59] & x[112]);
  assign t[203] = (x[95] & x[114]);
  assign t[204] = (x[95] & x[116]);
  assign t[205] = (x[88] & x[118]);
  assign t[206] = (x[95] & x[120]);
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[120]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[43] & t[44]);
  assign t[28] = ~(t[45] & t[122]);
  assign t[29] = t[15] ? x[24] : x[23];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[31];
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[39];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = ~(t[56] & t[123]);
  assign t[37] = t[15] ? x[29] : x[28];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[61] ^ t[62];
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[124]);
  assign t[44] = ~(t[125]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[71] & t[126]);
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = ~(t[74] & t[127]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[75] ? x[41] : x[40];
  assign t[51] = ~(t[76] & t[77]);
  assign t[52] = ~(t[78] & t[128]);
  assign t[53] = t[75] ? x[46] : x[45];
  assign t[54] = ~(t[129]);
  assign t[55] = ~(t[130]);
  assign t[56] = ~(t[79] & t[80]);
  assign t[57] = ~(t[81] & t[82]);
  assign t[58] = ~(t[83] & t[131]);
  assign t[59] = ~(t[84] & t[85]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[86] & t[132]);
  assign t[61] = t[87] ? x[58] : x[57];
  assign t[62] = ~(t[88] & t[89]);
  assign t[63] = ~(t[90] & t[91]);
  assign t[64] = ~(t[92] & t[133]);
  assign t[65] = t[87] ? x[63] : x[62];
  assign t[66] = ~(t[93] & t[94]);
  assign t[67] = ~(t[125] & t[124]);
  assign t[68] = ~(t[134]);
  assign t[69] = ~(t[135]);
  assign t[6] = ~(t[118] & t[119]);
  assign t[70] = ~(t[136]);
  assign t[71] = ~(t[95] & t[96]);
  assign t[72] = ~(t[137]);
  assign t[73] = ~(t[138]);
  assign t[74] = ~(t[97] & t[98]);
  assign t[75] = ~(t[22]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[130] & t[129]);
  assign t[7] = ~(t[120] & t[121]);
  assign t[80] = ~(t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[101] & t[102]);
  assign t[84] = ~(t[144]);
  assign t[85] = ~(t[145]);
  assign t[86] = ~(t[103] & t[104]);
  assign t[87] = ~(t[22]);
  assign t[88] = ~(t[105] & t[106]);
  assign t[89] = ~(t[107] & t[146]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[147]);
  assign t[91] = ~(t[148]);
  assign t[92] = ~(t[108] & t[109]);
  assign t[93] = ~(t[110] & t[111]);
  assign t[94] = ~(t[112] & t[149]);
  assign t[95] = ~(t[136] & t[135]);
  assign t[96] = ~(t[150]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[151]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[117];
endmodule

module R1ind152(x, y);
 input [101:0] x;
 output y;

 wire [166:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[135] ^ x[14];
  assign t[101] = t[136] ^ x[17];
  assign t[102] = t[137] ^ x[22];
  assign t[103] = t[138] ^ x[24];
  assign t[104] = t[139] ^ x[29];
  assign t[105] = t[140] ^ x[31];
  assign t[106] = t[141] ^ x[35];
  assign t[107] = t[142] ^ x[38];
  assign t[108] = t[143] ^ x[40];
  assign t[109] = t[144] ^ x[43];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[145] ^ x[45];
  assign t[111] = t[146] ^ x[50];
  assign t[112] = t[147] ^ x[52];
  assign t[113] = t[148] ^ x[56];
  assign t[114] = t[149] ^ x[59];
  assign t[115] = t[150] ^ x[61];
  assign t[116] = t[151] ^ x[64];
  assign t[117] = t[152] ^ x[66];
  assign t[118] = t[153] ^ x[71];
  assign t[119] = t[154] ^ x[73];
  assign t[11] = t[15] ? x[19] : x[18];
  assign t[120] = t[155] ^ x[77];
  assign t[121] = t[156] ^ x[79];
  assign t[122] = t[157] ^ x[81];
  assign t[123] = t[158] ^ x[83];
  assign t[124] = t[159] ^ x[85];
  assign t[125] = t[160] ^ x[88];
  assign t[126] = t[161] ^ x[90];
  assign t[127] = t[162] ^ x[92];
  assign t[128] = t[163] ^ x[95];
  assign t[129] = t[164] ^ x[97];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[165] ^ x[99];
  assign t[131] = t[166] ^ x[101];
  assign t[132] = (x[0] & x[1]);
  assign t[133] = (x[6] & x[7]);
  assign t[134] = (x[9] & x[10]);
  assign t[135] = (x[12] & x[13]);
  assign t[136] = (x[15] & x[16]);
  assign t[137] = (x[20] & x[21]);
  assign t[138] = (x[20] & x[23]);
  assign t[139] = (x[27] & x[28]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (x[27] & x[30]);
  assign t[141] = (x[20] & x[34]);
  assign t[142] = (x[36] & x[37]);
  assign t[143] = (x[36] & x[39]);
  assign t[144] = (x[41] & x[42]);
  assign t[145] = (x[41] & x[44]);
  assign t[146] = (x[48] & x[49]);
  assign t[147] = (x[48] & x[51]);
  assign t[148] = (x[27] & x[55]);
  assign t[149] = (x[57] & x[58]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (x[57] & x[60]);
  assign t[151] = (x[62] & x[63]);
  assign t[152] = (x[62] & x[65]);
  assign t[153] = (x[69] & x[70]);
  assign t[154] = (x[69] & x[72]);
  assign t[155] = (x[36] & x[76]);
  assign t[156] = (x[41] & x[78]);
  assign t[157] = (x[48] & x[80]);
  assign t[158] = (x[57] & x[82]);
  assign t[159] = (x[62] & x[84]);
  assign t[15] = ~(t[22]);
  assign t[160] = (x[86] & x[87]);
  assign t[161] = (x[86] & x[89]);
  assign t[162] = (x[69] & x[91]);
  assign t[163] = (x[93] & x[94]);
  assign t[164] = (x[93] & x[96]);
  assign t[165] = (x[86] & x[98]);
  assign t[166] = (x[93] & x[100]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[100]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[102] & t[43]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[29] = t[15] ? x[26] : x[25];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[31] = ~(t[47] & t[48]);
  assign t[32] = t[49] ^ t[39];
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[33];
  assign t[35] = ~(t[104] & t[53]);
  assign t[36] = ~(t[105] & t[54]);
  assign t[37] = t[15] ? x[33] : x[32];
  assign t[38] = ~(t[55] & t[56]);
  assign t[39] = ~(t[57] & t[58]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[59] ^ t[60];
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[106]);
  assign t[44] = ~(t[106] & t[65]);
  assign t[45] = ~(t[107] & t[66]);
  assign t[46] = ~(t[108] & t[67]);
  assign t[47] = ~(t[109] & t[68]);
  assign t[48] = ~(t[110] & t[69]);
  assign t[49] = t[70] ? x[47] : x[46];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = t[70] ? x[54] : x[53];
  assign t[53] = ~(t[113]);
  assign t[54] = ~(t[113] & t[73]);
  assign t[55] = ~(t[114] & t[74]);
  assign t[56] = ~(t[115] & t[75]);
  assign t[57] = ~(t[116] & t[76]);
  assign t[58] = ~(t[117] & t[77]);
  assign t[59] = t[78] ? x[68] : x[67];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[79] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = t[78] ? x[75] : x[74];
  assign t[64] = ~(t[83] & t[84]);
  assign t[65] = ~(t[102]);
  assign t[66] = ~(t[120]);
  assign t[67] = ~(t[120] & t[85]);
  assign t[68] = ~(t[121]);
  assign t[69] = ~(t[121] & t[86]);
  assign t[6] = ~(t[98] & t[99]);
  assign t[70] = ~(t[22]);
  assign t[71] = ~(t[122]);
  assign t[72] = ~(t[122] & t[87]);
  assign t[73] = ~(t[104]);
  assign t[74] = ~(t[123]);
  assign t[75] = ~(t[123] & t[88]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[124] & t[89]);
  assign t[78] = ~(t[22]);
  assign t[79] = ~(t[125] & t[90]);
  assign t[7] = ~(t[100] & t[101]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[127] & t[92]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[107]);
  assign t[86] = ~(t[109]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[114]);
  assign t[89] = ~(t[116]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[130]);
  assign t[91] = ~(t[130] & t[95]);
  assign t[92] = ~(t[118]);
  assign t[93] = ~(t[131]);
  assign t[94] = ~(t[131] & t[96]);
  assign t[95] = ~(t[125]);
  assign t[96] = ~(t[128]);
  assign t[97] = t[132] ^ x[2];
  assign t[98] = t[133] ^ x[8];
  assign t[99] = t[134] ^ x[11];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[97];
endmodule

module R1ind153(x, y);
 input [121:0] x;
 output y;

 wire [289:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[138] & t[139]);
  assign t[101] = ~(t[224]);
  assign t[102] = ~(t[212] | t[213]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[226]);
  assign t[105] = ~(t[140] | t[141]);
  assign t[106] = ~(t[138] & t[142]);
  assign t[107] = ~(t[227]);
  assign t[108] = ~(t[228]);
  assign t[109] = ~(t[143] | t[144]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[145] | t[146]);
  assign t[111] = ~(t[229] | t[147]);
  assign t[112] = t[148] ? x[88] : x[87];
  assign t[113] = ~(t[149] & t[150]);
  assign t[114] = ~(t[230]);
  assign t[115] = ~(t[231]);
  assign t[116] = ~(t[151] | t[152]);
  assign t[117] = ~(t[153] | t[154]);
  assign t[118] = ~(t[232] | t[155]);
  assign t[119] = t[148] ? x[97] : x[96];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[156] & t[142]);
  assign t[121] = ~(t[203]);
  assign t[122] = ~(t[157] & t[158]);
  assign t[123] = ~(t[159] & t[204]);
  assign t[124] = ~(t[80] | t[160]);
  assign t[125] = ~(t[80] | t[161]);
  assign t[126] = ~(x[4] & t[162]);
  assign t[127] = ~(t[204] & t[163]);
  assign t[128] = ~(t[233]);
  assign t[129] = ~(t[218] | t[219]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[156] & t[138]);
  assign t[131] = ~(t[80] | t[164]);
  assign t[132] = ~(t[234]);
  assign t[133] = ~(t[220] | t[221]);
  assign t[134] = ~(t[48]);
  assign t[135] = ~(t[165] | t[166]);
  assign t[136] = ~(t[235]);
  assign t[137] = ~(t[222] | t[223]);
  assign t[138] = ~(t[167] | t[166]);
  assign t[139] = ~(t[168] | t[169]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[236]);
  assign t[141] = ~(t[225] | t[226]);
  assign t[142] = ~(t[170] & t[171]);
  assign t[143] = ~(t[237]);
  assign t[144] = ~(t[227] | t[228]);
  assign t[145] = ~(t[238]);
  assign t[146] = ~(t[239]);
  assign t[147] = ~(t[172] | t[173]);
  assign t[148] = ~(t[48]);
  assign t[149] = ~(t[174] | t[175]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[176] & t[177]);
  assign t[151] = ~(t[240]);
  assign t[152] = ~(t[230] | t[231]);
  assign t[153] = ~(t[241]);
  assign t[154] = ~(t[242]);
  assign t[155] = ~(t[178] | t[179]);
  assign t[156] = ~(t[49] | t[168]);
  assign t[157] = ~(x[4] | t[202]);
  assign t[158] = ~(t[204]);
  assign t[159] = x[4] & t[202];
  assign t[15] = ~(t[201] & t[202]);
  assign t[160] = t[201] ? t[181] : t[180];
  assign t[161] = t[201] ? t[183] : t[182];
  assign t[162] = ~(t[202] | t[204]);
  assign t[163] = ~(x[4] | t[184]);
  assign t[164] = t[201] ? t[122] : t[123];
  assign t[165] = ~(t[121] | t[185]);
  assign t[166] = ~(t[121] | t[186]);
  assign t[167] = ~(t[121] | t[187]);
  assign t[168] = ~(t[188] & t[189]);
  assign t[169] = ~(t[150] & t[190]);
  assign t[16] = ~(t[203] & t[204]);
  assign t[170] = ~(t[202] | t[158]);
  assign t[171] = t[80] & t[201];
  assign t[172] = ~(t[243]);
  assign t[173] = ~(t[238] | t[239]);
  assign t[174] = ~(t[191] & t[142]);
  assign t[175] = t[51] | t[192];
  assign t[176] = t[204] & t[193];
  assign t[177] = t[157] | t[159];
  assign t[178] = ~(t[244]);
  assign t[179] = ~(t[241] | t[242]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[163] & t[158]);
  assign t[181] = ~(x[4] & t[170]);
  assign t[182] = ~(t[157] & t[204]);
  assign t[183] = ~(t[159] & t[158]);
  assign t[184] = ~(t[202]);
  assign t[185] = t[201] ? t[122] : t[183];
  assign t[186] = t[201] ? t[180] : t[126];
  assign t[187] = t[201] ? t[183] : t[122];
  assign t[188] = ~(t[165] | t[194]);
  assign t[189] = ~(t[121] & t[195]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[121] | t[196];
  assign t[191] = ~(t[193] & t[197]);
  assign t[192] = ~(t[80] | t[198]);
  assign t[193] = ~(t[121] | t[201]);
  assign t[194] = ~(t[80] | t[199]);
  assign t[195] = ~(t[126] & t[127]);
  assign t[196] = t[201] ? t[126] : t[180];
  assign t[197] = ~(t[127] & t[181]);
  assign t[198] = t[201] ? t[182] : t[183];
  assign t[199] = t[201] ? t[180] : t[181];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[245] ^ x[2];
  assign t[201] = t[246] ^ x[10];
  assign t[202] = t[247] ^ x[13];
  assign t[203] = t[248] ^ x[16];
  assign t[204] = t[249] ^ x[19];
  assign t[205] = t[250] ^ x[22];
  assign t[206] = t[251] ^ x[25];
  assign t[207] = t[252] ^ x[27];
  assign t[208] = t[253] ^ x[29];
  assign t[209] = t[254] ^ x[32];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[255] ^ x[37];
  assign t[211] = t[256] ^ x[40];
  assign t[212] = t[257] ^ x[42];
  assign t[213] = t[258] ^ x[44];
  assign t[214] = t[259] ^ x[47];
  assign t[215] = t[260] ^ x[52];
  assign t[216] = t[261] ^ x[55];
  assign t[217] = t[262] ^ x[57];
  assign t[218] = t[263] ^ x[59];
  assign t[219] = t[264] ^ x[61];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[63];
  assign t[221] = t[266] ^ x[65];
  assign t[222] = t[267] ^ x[69];
  assign t[223] = t[268] ^ x[71];
  assign t[224] = t[269] ^ x[75];
  assign t[225] = t[270] ^ x[77];
  assign t[226] = t[271] ^ x[79];
  assign t[227] = t[272] ^ x[81];
  assign t[228] = t[273] ^ x[83];
  assign t[229] = t[274] ^ x[86];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[90];
  assign t[231] = t[276] ^ x[92];
  assign t[232] = t[277] ^ x[95];
  assign t[233] = t[278] ^ x[99];
  assign t[234] = t[279] ^ x[101];
  assign t[235] = t[280] ^ x[103];
  assign t[236] = t[281] ^ x[105];
  assign t[237] = t[282] ^ x[107];
  assign t[238] = t[283] ^ x[109];
  assign t[239] = t[284] ^ x[111];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[113];
  assign t[241] = t[286] ^ x[115];
  assign t[242] = t[287] ^ x[117];
  assign t[243] = t[288] ^ x[119];
  assign t[244] = t[289] ^ x[121];
  assign t[245] = (x[0] & x[1]);
  assign t[246] = (x[8] & x[9]);
  assign t[247] = (x[11] & x[12]);
  assign t[248] = (x[14] & x[15]);
  assign t[249] = (x[17] & x[18]);
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = (x[20] & x[21]);
  assign t[251] = (x[23] & x[24]);
  assign t[252] = (x[20] & x[26]);
  assign t[253] = (x[20] & x[28]);
  assign t[254] = (x[30] & x[31]);
  assign t[255] = (x[35] & x[36]);
  assign t[256] = (x[38] & x[39]);
  assign t[257] = (x[23] & x[41]);
  assign t[258] = (x[23] & x[43]);
  assign t[259] = (x[45] & x[46]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[50] & x[51]);
  assign t[261] = (x[53] & x[54]);
  assign t[262] = (x[20] & x[56]);
  assign t[263] = (x[30] & x[58]);
  assign t[264] = (x[30] & x[60]);
  assign t[265] = (x[35] & x[62]);
  assign t[266] = (x[35] & x[64]);
  assign t[267] = (x[38] & x[68]);
  assign t[268] = (x[38] & x[70]);
  assign t[269] = (x[23] & x[74]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[45] & x[76]);
  assign t[271] = (x[45] & x[78]);
  assign t[272] = (x[50] & x[80]);
  assign t[273] = (x[50] & x[82]);
  assign t[274] = (x[84] & x[85]);
  assign t[275] = (x[53] & x[89]);
  assign t[276] = (x[53] & x[91]);
  assign t[277] = (x[93] & x[94]);
  assign t[278] = (x[30] & x[98]);
  assign t[279] = (x[35] & x[100]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[38] & x[102]);
  assign t[281] = (x[45] & x[104]);
  assign t[282] = (x[50] & x[106]);
  assign t[283] = (x[84] & x[108]);
  assign t[284] = (x[84] & x[110]);
  assign t[285] = (x[53] & x[112]);
  assign t[286] = (x[93] & x[114]);
  assign t[287] = (x[93] & x[116]);
  assign t[288] = (x[84] & x[118]);
  assign t[289] = (x[93] & x[120]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[205] | t[54]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[36] = ~(t[59] | t[60]);
  assign t[37] = ~(t[36] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[46] ^ t[64]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[65] | t[66]);
  assign t[41] = ~(t[206] | t[67]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[47] = ~(t[78] ^ t[79]);
  assign t[48] = ~(t[203]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[82]);
  assign t[51] = ~(t[80] | t[83]);
  assign t[52] = ~(t[207]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[84] | t[85]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = ~(t[209] | t[88]);
  assign t[57] = t[29] ? x[34] : x[33];
  assign t[58] = ~(t[89] & t[90]);
  assign t[59] = ~(t[91] | t[92]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[210] | t[93]);
  assign t[61] = ~(t[94] ^ t[95]);
  assign t[62] = ~(t[96] | t[97]);
  assign t[63] = ~(t[211] | t[98]);
  assign t[64] = ~(t[99] ^ t[100]);
  assign t[65] = ~(t[212]);
  assign t[66] = ~(t[213]);
  assign t[67] = ~(t[101] | t[102]);
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = ~(t[214] | t[105]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[29] ? x[49] : x[48];
  assign t[71] = t[106] | t[51];
  assign t[72] = ~(t[107] | t[108]);
  assign t[73] = ~(t[215] | t[109]);
  assign t[74] = ~(t[110] | t[111]);
  assign t[75] = ~(t[112] ^ t[113]);
  assign t[76] = ~(t[114] | t[115]);
  assign t[77] = ~(t[216] | t[116]);
  assign t[78] = ~(t[117] | t[118]);
  assign t[79] = ~(t[119] ^ t[120]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121]);
  assign t[81] = t[201] ? t[123] : t[122];
  assign t[82] = ~(t[124] | t[125]);
  assign t[83] = t[201] ? t[127] : t[126];
  assign t[84] = ~(t[217]);
  assign t[85] = ~(t[207] | t[208]);
  assign t[86] = ~(t[218]);
  assign t[87] = ~(t[219]);
  assign t[88] = ~(t[128] | t[129]);
  assign t[89] = ~(t[124] | t[130]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[131]);
  assign t[91] = ~(t[220]);
  assign t[92] = ~(t[221]);
  assign t[93] = ~(t[132] | t[133]);
  assign t[94] = t[134] ? x[67] : x[66];
  assign t[95] = ~(t[135] & t[31]);
  assign t[96] = ~(t[222]);
  assign t[97] = ~(t[223]);
  assign t[98] = ~(t[136] | t[137]);
  assign t[99] = t[134] ? x[73] : x[72];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[200];
endmodule

module R1ind154(x, y);
 input [121:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[108] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[31];
  assign t[117] = t[162] ^ x[33];
  assign t[118] = t[163] ^ x[36];
  assign t[119] = t[164] ^ x[39];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[44];
  assign t[121] = t[166] ^ x[48];
  assign t[122] = t[167] ^ x[50];
  assign t[123] = t[168] ^ x[53];
  assign t[124] = t[169] ^ x[56];
  assign t[125] = t[170] ^ x[61];
  assign t[126] = t[171] ^ x[65];
  assign t[127] = t[172] ^ x[67];
  assign t[128] = t[173] ^ x[69];
  assign t[129] = t[174] ^ x[71];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[73];
  assign t[131] = t[176] ^ x[76];
  assign t[132] = t[177] ^ x[78];
  assign t[133] = t[178] ^ x[80];
  assign t[134] = t[179] ^ x[82];
  assign t[135] = t[180] ^ x[84];
  assign t[136] = t[181] ^ x[86];
  assign t[137] = t[182] ^ x[88];
  assign t[138] = t[183] ^ x[90];
  assign t[139] = t[184] ^ x[92];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[94];
  assign t[141] = t[186] ^ x[97];
  assign t[142] = t[187] ^ x[99];
  assign t[143] = t[188] ^ x[101];
  assign t[144] = t[189] ^ x[103];
  assign t[145] = t[190] ^ x[105];
  assign t[146] = t[191] ^ x[107];
  assign t[147] = t[192] ^ x[109];
  assign t[148] = t[193] ^ x[111];
  assign t[149] = t[194] ^ x[113];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[115];
  assign t[151] = t[196] ^ x[117];
  assign t[152] = t[197] ^ x[119];
  assign t[153] = t[198] ^ x[121];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[20] & x[30]);
  assign t[162] = (x[20] & x[32]);
  assign t[163] = (x[34] & x[35]);
  assign t[164] = (x[37] & x[38]);
  assign t[165] = (x[42] & x[43]);
  assign t[166] = (x[25] & x[47]);
  assign t[167] = (x[25] & x[49]);
  assign t[168] = (x[51] & x[52]);
  assign t[169] = (x[54] & x[55]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[59] & x[60]);
  assign t[171] = (x[20] & x[64]);
  assign t[172] = (x[34] & x[66]);
  assign t[173] = (x[34] & x[68]);
  assign t[174] = (x[37] & x[70]);
  assign t[175] = (x[37] & x[72]);
  assign t[176] = (x[74] & x[75]);
  assign t[177] = (x[42] & x[77]);
  assign t[178] = (x[42] & x[79]);
  assign t[179] = (x[25] & x[81]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[51] & x[83]);
  assign t[181] = (x[51] & x[85]);
  assign t[182] = (x[54] & x[87]);
  assign t[183] = (x[54] & x[89]);
  assign t[184] = (x[59] & x[91]);
  assign t[185] = (x[59] & x[93]);
  assign t[186] = (x[95] & x[96]);
  assign t[187] = (x[34] & x[98]);
  assign t[188] = (x[37] & x[100]);
  assign t[189] = (x[74] & x[102]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[74] & x[104]);
  assign t[191] = (x[42] & x[106]);
  assign t[192] = (x[51] & x[108]);
  assign t[193] = (x[54] & x[110]);
  assign t[194] = (x[59] & x[112]);
  assign t[195] = (x[95] & x[114]);
  assign t[196] = (x[95] & x[116]);
  assign t[197] = (x[74] & x[118]);
  assign t[198] = (x[95] & x[120]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] ^ t[33];
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = t[60] | t[115];
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[43];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[69];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[70] | t[45]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[73] | t[118];
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = t[76] | t[119];
  assign t[53] = t[17] ? x[41] : x[40];
  assign t[54] = ~(t[77] & t[78]);
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = t[81] | t[120];
  assign t[57] = t[17] ? x[46] : x[45];
  assign t[58] = ~(t[121]);
  assign t[59] = ~(t[122]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[82] | t[58]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = t[85] | t[123];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = t[88] | t[124];
  assign t[65] = t[89] ? x[58] : x[57];
  assign t[66] = ~(t[90] & t[91]);
  assign t[67] = t[92] | t[125];
  assign t[68] = t[89] ? x[63] : x[62];
  assign t[69] = ~(t[93] & t[94]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[95] | t[71]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[96] | t[74]);
  assign t[77] = ~(t[97] & t[98]);
  assign t[78] = t[99] | t[131];
  assign t[79] = ~(t[132]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[100] | t[79]);
  assign t[82] = ~(t[134]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[101] | t[83]);
  assign t[86] = ~(t[137]);
  assign t[87] = ~(t[138]);
  assign t[88] = ~(t[102] | t[86]);
  assign t[89] = ~(t[24]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[139]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[103] | t[90]);
  assign t[93] = ~(t[104] & t[105]);
  assign t[94] = t[106] | t[141];
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[107] | t[97]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind155(x, y);
 input [121:0] x;
 output y;

 wire [207:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[114] & t[115]);
  assign t[103] = ~(t[142] & t[141]);
  assign t[104] = ~(t[155]);
  assign t[105] = ~(t[145] & t[144]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[147] & t[146]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[116] & t[117]);
  assign t[114] = ~(t[154] & t[153]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[160] & t[159]);
  assign t[117] = ~(t[162]);
  assign t[118] = t[163] ^ x[2];
  assign t[119] = t[164] ^ x[10];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[165] ^ x[13];
  assign t[121] = t[166] ^ x[16];
  assign t[122] = t[167] ^ x[19];
  assign t[123] = t[168] ^ x[22];
  assign t[124] = t[169] ^ x[27];
  assign t[125] = t[170] ^ x[31];
  assign t[126] = t[171] ^ x[33];
  assign t[127] = t[172] ^ x[36];
  assign t[128] = t[173] ^ x[39];
  assign t[129] = t[174] ^ x[44];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[48];
  assign t[131] = t[176] ^ x[50];
  assign t[132] = t[177] ^ x[53];
  assign t[133] = t[178] ^ x[56];
  assign t[134] = t[179] ^ x[61];
  assign t[135] = t[180] ^ x[65];
  assign t[136] = t[181] ^ x[67];
  assign t[137] = t[182] ^ x[69];
  assign t[138] = t[183] ^ x[71];
  assign t[139] = t[184] ^ x[73];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[76];
  assign t[141] = t[186] ^ x[78];
  assign t[142] = t[187] ^ x[80];
  assign t[143] = t[188] ^ x[82];
  assign t[144] = t[189] ^ x[84];
  assign t[145] = t[190] ^ x[86];
  assign t[146] = t[191] ^ x[88];
  assign t[147] = t[192] ^ x[90];
  assign t[148] = t[193] ^ x[92];
  assign t[149] = t[194] ^ x[94];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[97];
  assign t[151] = t[196] ^ x[99];
  assign t[152] = t[197] ^ x[101];
  assign t[153] = t[198] ^ x[103];
  assign t[154] = t[199] ^ x[105];
  assign t[155] = t[200] ^ x[107];
  assign t[156] = t[201] ^ x[109];
  assign t[157] = t[202] ^ x[111];
  assign t[158] = t[203] ^ x[113];
  assign t[159] = t[204] ^ x[115];
  assign t[15] = ~(t[119] & t[120]);
  assign t[160] = t[205] ^ x[117];
  assign t[161] = t[206] ^ x[119];
  assign t[162] = t[207] ^ x[121];
  assign t[163] = (x[0] & x[1]);
  assign t[164] = (x[8] & x[9]);
  assign t[165] = (x[11] & x[12]);
  assign t[166] = (x[14] & x[15]);
  assign t[167] = (x[17] & x[18]);
  assign t[168] = (x[20] & x[21]);
  assign t[169] = (x[25] & x[26]);
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = (x[20] & x[30]);
  assign t[171] = (x[20] & x[32]);
  assign t[172] = (x[34] & x[35]);
  assign t[173] = (x[37] & x[38]);
  assign t[174] = (x[42] & x[43]);
  assign t[175] = (x[25] & x[47]);
  assign t[176] = (x[25] & x[49]);
  assign t[177] = (x[51] & x[52]);
  assign t[178] = (x[54] & x[55]);
  assign t[179] = (x[59] & x[60]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[20] & x[64]);
  assign t[181] = (x[34] & x[66]);
  assign t[182] = (x[34] & x[68]);
  assign t[183] = (x[37] & x[70]);
  assign t[184] = (x[37] & x[72]);
  assign t[185] = (x[74] & x[75]);
  assign t[186] = (x[42] & x[77]);
  assign t[187] = (x[42] & x[79]);
  assign t[188] = (x[25] & x[81]);
  assign t[189] = (x[51] & x[83]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[51] & x[85]);
  assign t[191] = (x[54] & x[87]);
  assign t[192] = (x[54] & x[89]);
  assign t[193] = (x[59] & x[91]);
  assign t[194] = (x[59] & x[93]);
  assign t[195] = (x[95] & x[96]);
  assign t[196] = (x[34] & x[98]);
  assign t[197] = (x[37] & x[100]);
  assign t[198] = (x[74] & x[102]);
  assign t[199] = (x[74] & x[104]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[42] & x[106]);
  assign t[201] = (x[51] & x[108]);
  assign t[202] = (x[54] & x[110]);
  assign t[203] = (x[59] & x[112]);
  assign t[204] = (x[95] & x[114]);
  assign t[205] = (x[95] & x[116]);
  assign t[206] = (x[74] & x[118]);
  assign t[207] = (x[95] & x[120]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[121]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] & t[123]);
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] ^ t[33];
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = ~(t[60] & t[124]);
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[43];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[69];
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[74] & t[127]);
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = ~(t[77] & t[128]);
  assign t[53] = t[17] ? x[41] : x[40];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[80] & t[81]);
  assign t[56] = ~(t[82] & t[129]);
  assign t[57] = t[121] ? x[46] : x[45];
  assign t[58] = ~(t[130]);
  assign t[59] = ~(t[131]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[87] & t[132]);
  assign t[63] = ~(t[88] & t[89]);
  assign t[64] = ~(t[90] & t[133]);
  assign t[65] = t[48] ? x[58] : x[57];
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = ~(t[93] & t[134]);
  assign t[68] = t[48] ? x[63] : x[62];
  assign t[69] = ~(t[94] & t[95]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126] & t[125]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[96] & t[97]);
  assign t[75] = ~(t[138]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[98] & t[99]);
  assign t[78] = ~(t[100] & t[101]);
  assign t[79] = ~(t[102] & t[140]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[103] & t[104]);
  assign t[83] = ~(t[131] & t[130]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[105] & t[106]);
  assign t[88] = ~(t[146]);
  assign t[89] = ~(t[147]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[107] & t[108]);
  assign t[91] = ~(t[148]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[109] & t[110]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[113] & t[150]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[118];
endmodule

module R1ind156(x, y);
 input [101:0] x;
 output y;

 wire [167:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[135] ^ x[13];
  assign t[101] = t[136] ^ x[16];
  assign t[102] = t[137] ^ x[19];
  assign t[103] = t[138] ^ x[22];
  assign t[104] = t[139] ^ x[24];
  assign t[105] = t[140] ^ x[29];
  assign t[106] = t[141] ^ x[31];
  assign t[107] = t[142] ^ x[35];
  assign t[108] = t[143] ^ x[38];
  assign t[109] = t[144] ^ x[40];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] ^ x[43];
  assign t[111] = t[146] ^ x[45];
  assign t[112] = t[147] ^ x[50];
  assign t[113] = t[148] ^ x[52];
  assign t[114] = t[149] ^ x[56];
  assign t[115] = t[150] ^ x[59];
  assign t[116] = t[151] ^ x[61];
  assign t[117] = t[152] ^ x[64];
  assign t[118] = t[153] ^ x[66];
  assign t[119] = t[154] ^ x[71];
  assign t[11] = t[17] ? x[7] : x[6];
  assign t[120] = t[155] ^ x[73];
  assign t[121] = t[156] ^ x[77];
  assign t[122] = t[157] ^ x[79];
  assign t[123] = t[158] ^ x[81];
  assign t[124] = t[159] ^ x[84];
  assign t[125] = t[160] ^ x[86];
  assign t[126] = t[161] ^ x[88];
  assign t[127] = t[162] ^ x[90];
  assign t[128] = t[163] ^ x[93];
  assign t[129] = t[164] ^ x[95];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[165] ^ x[97];
  assign t[131] = t[166] ^ x[99];
  assign t[132] = t[167] ^ x[101];
  assign t[133] = (x[0] & x[1]);
  assign t[134] = (x[8] & x[9]);
  assign t[135] = (x[11] & x[12]);
  assign t[136] = (x[14] & x[15]);
  assign t[137] = (x[17] & x[18]);
  assign t[138] = (x[20] & x[21]);
  assign t[139] = (x[20] & x[23]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[27] & x[28]);
  assign t[141] = (x[27] & x[30]);
  assign t[142] = (x[20] & x[34]);
  assign t[143] = (x[36] & x[37]);
  assign t[144] = (x[36] & x[39]);
  assign t[145] = (x[41] & x[42]);
  assign t[146] = (x[41] & x[44]);
  assign t[147] = (x[48] & x[49]);
  assign t[148] = (x[48] & x[51]);
  assign t[149] = (x[27] & x[55]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[57] & x[58]);
  assign t[151] = (x[57] & x[60]);
  assign t[152] = (x[62] & x[63]);
  assign t[153] = (x[62] & x[65]);
  assign t[154] = (x[69] & x[70]);
  assign t[155] = (x[69] & x[72]);
  assign t[156] = (x[36] & x[76]);
  assign t[157] = (x[41] & x[78]);
  assign t[158] = (x[48] & x[80]);
  assign t[159] = (x[82] & x[83]);
  assign t[15] = ~(t[99] & t[100]);
  assign t[160] = (x[82] & x[85]);
  assign t[161] = (x[57] & x[87]);
  assign t[162] = (x[62] & x[89]);
  assign t[163] = (x[91] & x[92]);
  assign t[164] = (x[91] & x[94]);
  assign t[165] = (x[69] & x[96]);
  assign t[166] = (x[82] & x[98]);
  assign t[167] = (x[91] & x[100]);
  assign t[16] = ~(t[101] & t[102]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[101]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[103] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[104] & t[46]);
  assign t[31] = t[17] ? x[26] : x[25];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = t[51] ^ t[35];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[55];
  assign t[37] = ~(t[105] & t[56]);
  assign t[38] = ~(t[106] & t[57]);
  assign t[39] = t[17] ? x[33] : x[32];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[41];
  assign t[45] = ~(t[107]);
  assign t[46] = ~(t[107] & t[67]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = t[72] ? x[47] : x[46];
  assign t[52] = ~(t[112] & t[73]);
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = t[17] ? x[54] : x[53];
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[114] & t[77]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = t[72] ? x[68] : x[67];
  assign t[63] = ~(t[82] & t[83]);
  assign t[64] = ~(t[119] & t[84]);
  assign t[65] = ~(t[120] & t[85]);
  assign t[66] = t[72] ? x[75] : x[74];
  assign t[67] = ~(t[103]);
  assign t[68] = ~(t[121]);
  assign t[69] = ~(t[121] & t[86]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[24]);
  assign t[73] = ~(t[123]);
  assign t[74] = ~(t[123] & t[88]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[105]);
  assign t[78] = ~(t[126]);
  assign t[79] = ~(t[126] & t[91]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[131]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[131] & t[96]);
  assign t[91] = ~(t[115]);
  assign t[92] = ~(t[117]);
  assign t[93] = ~(t[132]);
  assign t[94] = ~(t[132] & t[97]);
  assign t[95] = ~(t[119]);
  assign t[96] = ~(t[124]);
  assign t[97] = ~(t[128]);
  assign t[98] = t[133] ^ x[2];
  assign t[99] = t[134] ^ x[10];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[98];
endmodule

module R1ind157(x, y);
 input [121:0] x;
 output y;

 wire [294:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[29] ? x[70] : x[69];
  assign t[101] = ~(t[142] & t[143]);
  assign t[102] = ~(t[228]);
  assign t[103] = ~(t[229]);
  assign t[104] = ~(t[144] | t[145]);
  assign t[105] = t[29] ? x[76] : x[75];
  assign t[106] = ~(t[146] & t[147]);
  assign t[107] = ~(t[230]);
  assign t[108] = ~(t[217] | t[218]);
  assign t[109] = ~(t[231]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[232]);
  assign t[111] = ~(t[148] | t[149]);
  assign t[112] = ~(t[150] | t[151]);
  assign t[113] = ~(t[233]);
  assign t[114] = ~(t[234]);
  assign t[115] = ~(t[152] | t[153]);
  assign t[116] = t[154] ? x[88] : x[87];
  assign t[117] = t[155] | t[83];
  assign t[118] = ~(t[235]);
  assign t[119] = ~(t[236]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[156] | t[157]);
  assign t[121] = ~(t[158] | t[159]);
  assign t[122] = ~(t[237] | t[160]);
  assign t[123] = t[154] ? x[97] : x[96];
  assign t[124] = ~(t[161] & t[162]);
  assign t[125] = ~(t[163] & t[164]);
  assign t[126] = ~(t[207] | t[165]);
  assign t[127] = t[128] & t[206];
  assign t[128] = ~(t[131]);
  assign t[129] = t[206] ? t[163] : t[166];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = t[206] ? t[168] : t[167];
  assign t[131] = ~(t[208]);
  assign t[132] = ~(t[238]);
  assign t[133] = ~(t[223] | t[224]);
  assign t[134] = ~(t[131] | t[169]);
  assign t[135] = ~(t[128] | t[170]);
  assign t[136] = ~(t[171] & t[172]);
  assign t[137] = ~(t[239]);
  assign t[138] = ~(t[225] | t[226]);
  assign t[139] = ~(t[240]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[241]);
  assign t[141] = ~(t[173] | t[174]);
  assign t[142] = ~(t[150] | t[175]);
  assign t[143] = ~(t[117] | t[176]);
  assign t[144] = ~(t[242]);
  assign t[145] = ~(t[228] | t[229]);
  assign t[146] = ~(t[177] | t[84]);
  assign t[147] = ~(t[134] | t[155]);
  assign t[148] = ~(t[243]);
  assign t[149] = ~(t[231] | t[232]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[128] | t[178]);
  assign t[151] = ~(t[93] & t[179]);
  assign t[152] = ~(t[244]);
  assign t[153] = ~(t[233] | t[234]);
  assign t[154] = ~(t[48]);
  assign t[155] = ~(t[180] & t[82]);
  assign t[156] = ~(t[245]);
  assign t[157] = ~(t[235] | t[236]);
  assign t[158] = ~(t[246]);
  assign t[159] = ~(t[247]);
  assign t[15] = ~(t[206] & t[207]);
  assign t[160] = ~(t[181] | t[182]);
  assign t[161] = ~(t[150]);
  assign t[162] = ~(t[183] | t[83]);
  assign t[163] = ~(t[209] & t[184]);
  assign t[164] = ~(x[4] & t[126]);
  assign t[165] = ~(t[209]);
  assign t[166] = ~(x[4] & t[185]);
  assign t[167] = ~(t[87] & t[165]);
  assign t[168] = ~(t[86] & t[209]);
  assign t[169] = t[206] ? t[186] : t[167];
  assign t[16] = ~(t[208] & t[209]);
  assign t[170] = t[206] ? t[187] : t[164];
  assign t[171] = ~(t[150] | t[188]);
  assign t[172] = t[131] | t[189];
  assign t[173] = ~(t[248]);
  assign t[174] = ~(t[240] | t[241]);
  assign t[175] = ~(t[128] | t[190]);
  assign t[176] = ~(t[191] & t[172]);
  assign t[177] = ~(t[128] | t[192]);
  assign t[178] = t[206] ? t[193] : t[186];
  assign t[179] = ~(t[131] & t[194]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[195] | t[196]);
  assign t[181] = ~(t[249]);
  assign t[182] = ~(t[246] | t[247]);
  assign t[183] = ~(t[197]);
  assign t[184] = ~(x[4] | t[198]);
  assign t[185] = ~(t[207] | t[209]);
  assign t[186] = ~(t[86] & t[165]);
  assign t[187] = ~(t[184] & t[165]);
  assign t[188] = ~(t[128] | t[199]);
  assign t[189] = t[206] ? t[166] : t[187];
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[206] ? t[166] : t[163];
  assign t[191] = ~(t[200] | t[201]);
  assign t[192] = t[206] ? t[186] : t[193];
  assign t[193] = ~(t[87] & t[209]);
  assign t[194] = ~(t[166] & t[163]);
  assign t[195] = ~(t[131] | t[202]);
  assign t[196] = ~(t[131] | t[203]);
  assign t[197] = ~(t[201] | t[188]);
  assign t[198] = ~(t[207]);
  assign t[199] = t[206] ? t[167] : t[168];
  assign t[19] = t[29] ? x[7] : x[6];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = ~(t[81]);
  assign t[201] = ~(t[128] | t[204]);
  assign t[202] = t[206] ? t[167] : t[186];
  assign t[203] = t[206] ? t[187] : t[166];
  assign t[204] = t[206] ? t[164] : t[187];
  assign t[205] = t[250] ^ x[2];
  assign t[206] = t[251] ^ x[10];
  assign t[207] = t[252] ^ x[13];
  assign t[208] = t[253] ^ x[16];
  assign t[209] = t[254] ^ x[19];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[255] ^ x[22];
  assign t[211] = t[256] ^ x[25];
  assign t[212] = t[257] ^ x[27];
  assign t[213] = t[258] ^ x[29];
  assign t[214] = t[259] ^ x[32];
  assign t[215] = t[260] ^ x[37];
  assign t[216] = t[261] ^ x[40];
  assign t[217] = t[262] ^ x[42];
  assign t[218] = t[263] ^ x[44];
  assign t[219] = t[264] ^ x[47];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[52];
  assign t[221] = t[266] ^ x[55];
  assign t[222] = t[267] ^ x[57];
  assign t[223] = t[268] ^ x[59];
  assign t[224] = t[269] ^ x[61];
  assign t[225] = t[270] ^ x[63];
  assign t[226] = t[271] ^ x[65];
  assign t[227] = t[272] ^ x[68];
  assign t[228] = t[273] ^ x[72];
  assign t[229] = t[274] ^ x[74];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[78];
  assign t[231] = t[276] ^ x[80];
  assign t[232] = t[277] ^ x[82];
  assign t[233] = t[278] ^ x[84];
  assign t[234] = t[279] ^ x[86];
  assign t[235] = t[280] ^ x[90];
  assign t[236] = t[281] ^ x[92];
  assign t[237] = t[282] ^ x[95];
  assign t[238] = t[283] ^ x[99];
  assign t[239] = t[284] ^ x[101];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[103];
  assign t[241] = t[286] ^ x[105];
  assign t[242] = t[287] ^ x[107];
  assign t[243] = t[288] ^ x[109];
  assign t[244] = t[289] ^ x[111];
  assign t[245] = t[290] ^ x[113];
  assign t[246] = t[291] ^ x[115];
  assign t[247] = t[292] ^ x[117];
  assign t[248] = t[293] ^ x[119];
  assign t[249] = t[294] ^ x[121];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = (x[0] & x[1]);
  assign t[251] = (x[8] & x[9]);
  assign t[252] = (x[11] & x[12]);
  assign t[253] = (x[14] & x[15]);
  assign t[254] = (x[17] & x[18]);
  assign t[255] = (x[20] & x[21]);
  assign t[256] = (x[23] & x[24]);
  assign t[257] = (x[20] & x[26]);
  assign t[258] = (x[20] & x[28]);
  assign t[259] = (x[30] & x[31]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[35] & x[36]);
  assign t[261] = (x[38] & x[39]);
  assign t[262] = (x[23] & x[41]);
  assign t[263] = (x[23] & x[43]);
  assign t[264] = (x[45] & x[46]);
  assign t[265] = (x[50] & x[51]);
  assign t[266] = (x[53] & x[54]);
  assign t[267] = (x[20] & x[56]);
  assign t[268] = (x[30] & x[58]);
  assign t[269] = (x[30] & x[60]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[35] & x[62]);
  assign t[271] = (x[35] & x[64]);
  assign t[272] = (x[66] & x[67]);
  assign t[273] = (x[38] & x[71]);
  assign t[274] = (x[38] & x[73]);
  assign t[275] = (x[23] & x[77]);
  assign t[276] = (x[45] & x[79]);
  assign t[277] = (x[45] & x[81]);
  assign t[278] = (x[50] & x[83]);
  assign t[279] = (x[50] & x[85]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[53] & x[89]);
  assign t[281] = (x[53] & x[91]);
  assign t[282] = (x[93] & x[94]);
  assign t[283] = (x[30] & x[98]);
  assign t[284] = (x[35] & x[100]);
  assign t[285] = (x[66] & x[102]);
  assign t[286] = (x[66] & x[104]);
  assign t[287] = (x[38] & x[106]);
  assign t[288] = (x[45] & x[108]);
  assign t[289] = (x[50] & x[110]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[290] = (x[53] & x[112]);
  assign t[291] = (x[93] & x[114]);
  assign t[292] = (x[93] & x[116]);
  assign t[293] = (x[66] & x[118]);
  assign t[294] = (x[93] & x[120]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51] & t[52]);
  assign t[32] = ~(t[53] | t[54]);
  assign t[33] = ~(t[210] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[58] ^ t[59]);
  assign t[36] = ~(t[60] | t[61]);
  assign t[37] = ~(t[62] ^ t[63]);
  assign t[38] = ~(t[64] | t[65]);
  assign t[39] = ~(t[36] ^ t[66]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[67] | t[68]);
  assign t[41] = ~(t[211] | t[69]);
  assign t[42] = ~(t[70] | t[71]);
  assign t[43] = ~(t[72] ^ t[73]);
  assign t[44] = ~(t[74] | t[75]);
  assign t[45] = ~(t[46] ^ t[76]);
  assign t[46] = ~(t[77] | t[78]);
  assign t[47] = ~(t[79] ^ t[80]);
  assign t[48] = ~(t[208]);
  assign t[49] = ~(t[81] & t[82]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[83] | t[84];
  assign t[51] = t[209] & t[85];
  assign t[52] = t[86] | t[87];
  assign t[53] = ~(t[212]);
  assign t[54] = ~(t[213]);
  assign t[55] = ~(t[88] | t[89]);
  assign t[56] = ~(t[90] | t[91]);
  assign t[57] = ~(t[214] | t[92]);
  assign t[58] = t[29] ? x[34] : x[33];
  assign t[59] = ~(t[93] & t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[215] | t[97]);
  assign t[62] = ~(t[98] | t[99]);
  assign t[63] = ~(t[100] ^ t[101]);
  assign t[64] = ~(t[102] | t[103]);
  assign t[65] = ~(t[216] | t[104]);
  assign t[66] = ~(t[105] ^ t[106]);
  assign t[67] = ~(t[217]);
  assign t[68] = ~(t[218]);
  assign t[69] = ~(t[107] | t[108]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[109] | t[110]);
  assign t[71] = ~(t[219] | t[111]);
  assign t[72] = t[29] ? x[49] : x[48];
  assign t[73] = ~(t[112] & t[82]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[220] | t[115]);
  assign t[76] = ~(t[116] ^ t[117]);
  assign t[77] = ~(t[118] | t[119]);
  assign t[78] = ~(t[221] | t[120]);
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[123] ^ t[124]);
  assign t[81] = ~(t[85] & t[125]);
  assign t[82] = ~(t[126] & t[127]);
  assign t[83] = ~(t[128] | t[129]);
  assign t[84] = ~(t[128] | t[130]);
  assign t[85] = ~(t[131] | t[206]);
  assign t[86] = ~(x[4] | t[207]);
  assign t[87] = x[4] & t[207];
  assign t[88] = ~(t[222]);
  assign t[89] = ~(t[212] | t[213]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[223]);
  assign t[91] = ~(t[224]);
  assign t[92] = ~(t[132] | t[133]);
  assign t[93] = ~(t[134] | t[135]);
  assign t[94] = ~(t[84] | t[136]);
  assign t[95] = ~(t[225]);
  assign t[96] = ~(t[226]);
  assign t[97] = ~(t[137] | t[138]);
  assign t[98] = ~(t[139] | t[140]);
  assign t[99] = ~(t[227] | t[141]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[205];
endmodule

module R1ind158(x, y);
 input [112:0] x;
 output y;

 wire [182:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141]);
  assign t[101] = t[142] ^ x[2];
  assign t[102] = t[143] ^ x[10];
  assign t[103] = t[144] ^ x[13];
  assign t[104] = t[145] ^ x[16];
  assign t[105] = t[146] ^ x[19];
  assign t[106] = t[147] ^ x[22];
  assign t[107] = t[148] ^ x[27];
  assign t[108] = t[149] ^ x[31];
  assign t[109] = t[150] ^ x[33];
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[36];
  assign t[111] = t[152] ^ x[41];
  assign t[112] = t[153] ^ x[45];
  assign t[113] = t[154] ^ x[47];
  assign t[114] = t[155] ^ x[50];
  assign t[115] = t[156] ^ x[53];
  assign t[116] = t[157] ^ x[58];
  assign t[117] = t[158] ^ x[62];
  assign t[118] = t[159] ^ x[64];
  assign t[119] = t[160] ^ x[66];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[69];
  assign t[121] = t[162] ^ x[71];
  assign t[122] = t[163] ^ x[73];
  assign t[123] = t[164] ^ x[75];
  assign t[124] = t[165] ^ x[77];
  assign t[125] = t[166] ^ x[79];
  assign t[126] = t[167] ^ x[81];
  assign t[127] = t[168] ^ x[83];
  assign t[128] = t[169] ^ x[85];
  assign t[129] = t[170] ^ x[87];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[90];
  assign t[131] = t[172] ^ x[92];
  assign t[132] = t[173] ^ x[94];
  assign t[133] = t[174] ^ x[96];
  assign t[134] = t[175] ^ x[98];
  assign t[135] = t[176] ^ x[100];
  assign t[136] = t[177] ^ x[102];
  assign t[137] = t[178] ^ x[104];
  assign t[138] = t[179] ^ x[106];
  assign t[139] = t[180] ^ x[108];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[110];
  assign t[141] = t[182] ^ x[112];
  assign t[142] = (x[0] & x[1]);
  assign t[143] = (x[8] & x[9]);
  assign t[144] = (x[11] & x[12]);
  assign t[145] = (x[14] & x[15]);
  assign t[146] = (x[17] & x[18]);
  assign t[147] = (x[20] & x[21]);
  assign t[148] = (x[25] & x[26]);
  assign t[149] = (x[20] & x[30]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[20] & x[32]);
  assign t[151] = (x[34] & x[35]);
  assign t[152] = (x[39] & x[40]);
  assign t[153] = (x[25] & x[44]);
  assign t[154] = (x[25] & x[46]);
  assign t[155] = (x[48] & x[49]);
  assign t[156] = (x[51] & x[52]);
  assign t[157] = (x[56] & x[57]);
  assign t[158] = (x[20] & x[61]);
  assign t[159] = (x[34] & x[63]);
  assign t[15] = ~(t[102] & t[103]);
  assign t[160] = (x[34] & x[65]);
  assign t[161] = (x[67] & x[68]);
  assign t[162] = (x[39] & x[70]);
  assign t[163] = (x[39] & x[72]);
  assign t[164] = (x[25] & x[74]);
  assign t[165] = (x[48] & x[76]);
  assign t[166] = (x[48] & x[78]);
  assign t[167] = (x[51] & x[80]);
  assign t[168] = (x[51] & x[82]);
  assign t[169] = (x[56] & x[84]);
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = (x[56] & x[86]);
  assign t[171] = (x[88] & x[89]);
  assign t[172] = (x[34] & x[91]);
  assign t[173] = (x[67] & x[93]);
  assign t[174] = (x[67] & x[95]);
  assign t[175] = (x[39] & x[97]);
  assign t[176] = (x[48] & x[99]);
  assign t[177] = (x[51] & x[101]);
  assign t[178] = (x[56] & x[103]);
  assign t[179] = (x[88] & x[105]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[88] & x[107]);
  assign t[181] = (x[67] & x[109]);
  assign t[182] = (x[88] & x[111]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[104]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] | t[106];
  assign t[31] = t[104] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[50];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[40];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] | t[107];
  assign t[38] = t[17] ? x[29] : x[28];
  assign t[39] = ~(t[57] & t[58]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = t[61] ^ t[42];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[108]);
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[66] | t[44]);
  assign t[47] = ~(t[67] & t[68]);
  assign t[48] = t[69] | t[110];
  assign t[49] = t[104] ? x[38] : x[37];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[70] & t[71]);
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = t[74] | t[111];
  assign t[53] = t[75] ? x[43] : x[42];
  assign t[54] = ~(t[112]);
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[76] | t[54]);
  assign t[57] = ~(t[77] & t[78]);
  assign t[58] = t[79] | t[114];
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[82] | t[115];
  assign t[61] = t[75] ? x[55] : x[54];
  assign t[62] = ~(t[83] & t[84]);
  assign t[63] = t[85] | t[116];
  assign t[64] = t[75] ? x[60] : x[59];
  assign t[65] = ~(t[86] & t[87]);
  assign t[66] = ~(t[117]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[88] | t[67]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[89] & t[90]);
  assign t[71] = t[91] | t[120];
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[92] | t[72]);
  assign t[75] = ~(t[24]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[93] | t[77]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[94] | t[80]);
  assign t[83] = ~(t[128]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[95] | t[83]);
  assign t[86] = ~(t[96] & t[97]);
  assign t[87] = t[98] | t[130];
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[99] | t[89]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[100] | t[96]);
  assign t[99] = ~(t[140]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[101];
endmodule

module R1ind159(x, y);
 input [112:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[145]);
  assign t[101] = ~(t[138] & t[137]);
  assign t[102] = ~(t[146]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[108] & t[109]);
  assign t[106] = ~(t[142] & t[141]);
  assign t[107] = ~(t[149]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[150]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[2];
  assign t[111] = t[152] ^ x[10];
  assign t[112] = t[153] ^ x[13];
  assign t[113] = t[154] ^ x[16];
  assign t[114] = t[155] ^ x[19];
  assign t[115] = t[156] ^ x[22];
  assign t[116] = t[157] ^ x[27];
  assign t[117] = t[158] ^ x[31];
  assign t[118] = t[159] ^ x[33];
  assign t[119] = t[160] ^ x[36];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[41];
  assign t[121] = t[162] ^ x[45];
  assign t[122] = t[163] ^ x[47];
  assign t[123] = t[164] ^ x[50];
  assign t[124] = t[165] ^ x[53];
  assign t[125] = t[166] ^ x[58];
  assign t[126] = t[167] ^ x[62];
  assign t[127] = t[168] ^ x[64];
  assign t[128] = t[169] ^ x[66];
  assign t[129] = t[170] ^ x[69];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[71];
  assign t[131] = t[172] ^ x[73];
  assign t[132] = t[173] ^ x[75];
  assign t[133] = t[174] ^ x[77];
  assign t[134] = t[175] ^ x[79];
  assign t[135] = t[176] ^ x[81];
  assign t[136] = t[177] ^ x[83];
  assign t[137] = t[178] ^ x[85];
  assign t[138] = t[179] ^ x[87];
  assign t[139] = t[180] ^ x[90];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[92];
  assign t[141] = t[182] ^ x[94];
  assign t[142] = t[183] ^ x[96];
  assign t[143] = t[184] ^ x[98];
  assign t[144] = t[185] ^ x[100];
  assign t[145] = t[186] ^ x[102];
  assign t[146] = t[187] ^ x[104];
  assign t[147] = t[188] ^ x[106];
  assign t[148] = t[189] ^ x[108];
  assign t[149] = t[190] ^ x[110];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[191] ^ x[112];
  assign t[151] = (x[0] & x[1]);
  assign t[152] = (x[8] & x[9]);
  assign t[153] = (x[11] & x[12]);
  assign t[154] = (x[14] & x[15]);
  assign t[155] = (x[17] & x[18]);
  assign t[156] = (x[20] & x[21]);
  assign t[157] = (x[25] & x[26]);
  assign t[158] = (x[20] & x[30]);
  assign t[159] = (x[20] & x[32]);
  assign t[15] = ~(t[111] & t[112]);
  assign t[160] = (x[34] & x[35]);
  assign t[161] = (x[39] & x[40]);
  assign t[162] = (x[25] & x[44]);
  assign t[163] = (x[25] & x[46]);
  assign t[164] = (x[48] & x[49]);
  assign t[165] = (x[51] & x[52]);
  assign t[166] = (x[56] & x[57]);
  assign t[167] = (x[20] & x[61]);
  assign t[168] = (x[34] & x[63]);
  assign t[169] = (x[34] & x[65]);
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = (x[67] & x[68]);
  assign t[171] = (x[39] & x[70]);
  assign t[172] = (x[39] & x[72]);
  assign t[173] = (x[25] & x[74]);
  assign t[174] = (x[48] & x[76]);
  assign t[175] = (x[48] & x[78]);
  assign t[176] = (x[51] & x[80]);
  assign t[177] = (x[51] & x[82]);
  assign t[178] = (x[56] & x[84]);
  assign t[179] = (x[56] & x[86]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[88] & x[89]);
  assign t[181] = (x[34] & x[91]);
  assign t[182] = (x[67] & x[93]);
  assign t[183] = (x[67] & x[95]);
  assign t[184] = (x[39] & x[97]);
  assign t[185] = (x[48] & x[99]);
  assign t[186] = (x[51] & x[101]);
  assign t[187] = (x[56] & x[103]);
  assign t[188] = (x[88] & x[105]);
  assign t[189] = (x[88] & x[107]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[67] & x[109]);
  assign t[191] = (x[88] & x[111]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[113]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[115]);
  assign t[31] = t[113] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[50];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[40];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = ~(t[56] & t[116]);
  assign t[38] = t[17] ? x[29] : x[28];
  assign t[39] = ~(t[57] & t[58]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = t[61] ^ t[42];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[117]);
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[66] & t[67]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = ~(t[70] & t[119]);
  assign t[49] = t[113] ? x[38] : x[37];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[71] & t[72]);
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[120]);
  assign t[53] = t[17] ? x[43] : x[42];
  assign t[54] = ~(t[121]);
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = ~(t[80] & t[123]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[83] & t[124]);
  assign t[61] = t[84] ? x[55] : x[54];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = ~(t[87] & t[125]);
  assign t[64] = t[84] ? x[60] : x[59];
  assign t[65] = ~(t[88] & t[89]);
  assign t[66] = ~(t[118] & t[117]);
  assign t[67] = ~(t[126]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[128]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[90] & t[91]);
  assign t[71] = ~(t[92] & t[93]);
  assign t[72] = ~(t[94] & t[129]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[95] & t[96]);
  assign t[76] = ~(t[122] & t[121]);
  assign t[77] = ~(t[132]);
  assign t[78] = ~(t[133]);
  assign t[79] = ~(t[134]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[97] & t[98]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[99] & t[100]);
  assign t[84] = ~(t[24]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[101] & t[102]);
  assign t[88] = ~(t[103] & t[104]);
  assign t[89] = ~(t[105] & t[139]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[106] & t[107]);
  assign t[95] = ~(t[131] & t[130]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[134] & t[133]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[110];
endmodule

module R1ind160(x, y);
 input [94:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[29];
  assign t[101] = t[133] ^ x[31];
  assign t[102] = t[134] ^ x[35];
  assign t[103] = t[135] ^ x[38];
  assign t[104] = t[136] ^ x[40];
  assign t[105] = t[137] ^ x[45];
  assign t[106] = t[138] ^ x[47];
  assign t[107] = t[139] ^ x[51];
  assign t[108] = t[140] ^ x[54];
  assign t[109] = t[141] ^ x[56];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[59];
  assign t[111] = t[143] ^ x[61];
  assign t[112] = t[144] ^ x[66];
  assign t[113] = t[145] ^ x[68];
  assign t[114] = t[146] ^ x[72];
  assign t[115] = t[147] ^ x[75];
  assign t[116] = t[148] ^ x[77];
  assign t[117] = t[149] ^ x[79];
  assign t[118] = t[150] ^ x[81];
  assign t[119] = t[151] ^ x[83];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[152] ^ x[86];
  assign t[121] = t[153] ^ x[88];
  assign t[122] = t[154] ^ x[90];
  assign t[123] = t[155] ^ x[92];
  assign t[124] = t[156] ^ x[94];
  assign t[125] = (x[0] & x[1]);
  assign t[126] = (x[8] & x[9]);
  assign t[127] = (x[11] & x[12]);
  assign t[128] = (x[14] & x[15]);
  assign t[129] = (x[17] & x[18]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & x[21]);
  assign t[131] = (x[20] & x[23]);
  assign t[132] = (x[27] & x[28]);
  assign t[133] = (x[27] & x[30]);
  assign t[134] = (x[20] & x[34]);
  assign t[135] = (x[36] & x[37]);
  assign t[136] = (x[36] & x[39]);
  assign t[137] = (x[43] & x[44]);
  assign t[138] = (x[43] & x[46]);
  assign t[139] = (x[27] & x[50]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[52] & x[53]);
  assign t[141] = (x[52] & x[55]);
  assign t[142] = (x[57] & x[58]);
  assign t[143] = (x[57] & x[60]);
  assign t[144] = (x[64] & x[65]);
  assign t[145] = (x[64] & x[67]);
  assign t[146] = (x[36] & x[71]);
  assign t[147] = (x[73] & x[74]);
  assign t[148] = (x[73] & x[76]);
  assign t[149] = (x[43] & x[78]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[52] & x[80]);
  assign t[151] = (x[57] & x[82]);
  assign t[152] = (x[84] & x[85]);
  assign t[153] = (x[84] & x[87]);
  assign t[154] = (x[64] & x[89]);
  assign t[155] = (x[73] & x[91]);
  assign t[156] = (x[84] & x[93]);
  assign t[15] = ~(t[94] & t[95]);
  assign t[16] = ~(t[96] & t[97]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[96]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[98] & t[44]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = t[96] ? x[26] : x[25];
  assign t[32] = ~(t[46] & t[47]);
  assign t[33] = t[48] ^ t[49];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[42];
  assign t[36] = ~(t[100] & t[53]);
  assign t[37] = ~(t[101] & t[54]);
  assign t[38] = t[17] ? x[33] : x[32];
  assign t[39] = ~(t[55] & t[56]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = t[59] ^ t[60];
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[40];
  assign t[44] = ~(t[102]);
  assign t[45] = ~(t[102] & t[64]);
  assign t[46] = ~(t[103] & t[65]);
  assign t[47] = ~(t[104] & t[66]);
  assign t[48] = t[96] ? x[42] : x[41];
  assign t[49] = ~(t[67] & t[68]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = t[71] ? x[49] : x[48];
  assign t[53] = ~(t[107]);
  assign t[54] = ~(t[107] & t[72]);
  assign t[55] = ~(t[108] & t[73]);
  assign t[56] = ~(t[109] & t[74]);
  assign t[57] = ~(t[110] & t[75]);
  assign t[58] = ~(t[111] & t[76]);
  assign t[59] = t[77] ? x[63] : x[62];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[78] & t[79]);
  assign t[61] = ~(t[112] & t[80]);
  assign t[62] = ~(t[113] & t[81]);
  assign t[63] = t[77] ? x[70] : x[69];
  assign t[64] = ~(t[98]);
  assign t[65] = ~(t[114]);
  assign t[66] = ~(t[114] & t[82]);
  assign t[67] = ~(t[115] & t[83]);
  assign t[68] = ~(t[116] & t[84]);
  assign t[69] = ~(t[117]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[117] & t[85]);
  assign t[71] = ~(t[24]);
  assign t[72] = ~(t[100]);
  assign t[73] = ~(t[118]);
  assign t[74] = ~(t[118] & t[86]);
  assign t[75] = ~(t[119]);
  assign t[76] = ~(t[119] & t[87]);
  assign t[77] = ~(t[24]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121] & t[89]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[122]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[123]);
  assign t[84] = ~(t[123] & t[91]);
  assign t[85] = ~(t[105]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[124]);
  assign t[89] = ~(t[124] & t[92]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[115]);
  assign t[92] = ~(t[120]);
  assign t[93] = t[125] ^ x[2];
  assign t[94] = t[126] ^ x[10];
  assign t[95] = t[127] ^ x[13];
  assign t[96] = t[128] ^ x[16];
  assign t[97] = t[129] ^ x[19];
  assign t[98] = t[130] ^ x[22];
  assign t[99] = t[131] ^ x[24];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[93];
endmodule

module R1ind161(x, y);
 input [112:0] x;
 output y;

 wire [275:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[205] | t[206]);
  assign t[101] = ~(t[217]);
  assign t[102] = ~(t[218]);
  assign t[103] = ~(t[137] | t[138]);
  assign t[104] = ~(t[85] | t[139]);
  assign t[105] = ~(t[140] & t[141]);
  assign t[106] = ~(t[219]);
  assign t[107] = ~(t[220]);
  assign t[108] = ~(t[142] | t[143]);
  assign t[109] = t[144] ? x[81] : x[80];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] | t[146];
  assign t[111] = ~(t[221]);
  assign t[112] = ~(t[222]);
  assign t[113] = ~(t[147] | t[148]);
  assign t[114] = ~(t[149] | t[150]);
  assign t[115] = ~(t[223] | t[151]);
  assign t[116] = t[144] ? x[90] : x[89];
  assign t[117] = ~(t[152] & t[153]);
  assign t[118] = ~(t[197]);
  assign t[119] = ~(t[154] & t[82]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[155] & t[198]);
  assign t[121] = ~(t[118] | t[156]);
  assign t[122] = ~(t[78] | t[157]);
  assign t[123] = ~(t[158] & t[159]);
  assign t[124] = ~(t[160] & t[161]);
  assign t[125] = ~(t[162] | t[163]);
  assign t[126] = ~(t[164] | t[165]);
  assign t[127] = ~(t[224]);
  assign t[128] = ~(t[211] | t[212]);
  assign t[129] = ~(t[162] | t[166]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[167] | t[168]);
  assign t[131] = ~(t[225]);
  assign t[132] = ~(t[213] | t[214]);
  assign t[133] = ~(t[226]);
  assign t[134] = ~(t[227]);
  assign t[135] = ~(t[169] | t[170]);
  assign t[136] = ~(t[171] | t[165]);
  assign t[137] = ~(t[228]);
  assign t[138] = ~(t[217] | t[218]);
  assign t[139] = t[146] | t[163];
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = t[198] & t[160];
  assign t[141] = t[154] | t[155];
  assign t[142] = ~(t[229]);
  assign t[143] = ~(t[219] | t[220]);
  assign t[144] = ~(t[47]);
  assign t[145] = ~(t[172] & t[31]);
  assign t[146] = ~(t[78] | t[173]);
  assign t[147] = ~(t[230]);
  assign t[148] = ~(t[221] | t[222]);
  assign t[149] = ~(t[231]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[232]);
  assign t[151] = ~(t[174] | t[175]);
  assign t[152] = ~(t[48]);
  assign t[153] = ~(t[176] | t[146]);
  assign t[154] = ~(x[4] | t[196]);
  assign t[155] = x[4] & t[196];
  assign t[156] = t[195] ? t[119] : t[177];
  assign t[157] = t[195] ? t[179] : t[178];
  assign t[158] = ~(x[4] & t[180]);
  assign t[159] = ~(t[198] & t[181]);
  assign t[15] = ~(t[195] & t[196]);
  assign t[160] = ~(t[118] | t[195]);
  assign t[161] = ~(t[159] & t[178]);
  assign t[162] = ~(t[78] | t[182]);
  assign t[163] = ~(t[78] | t[183]);
  assign t[164] = ~(t[78] | t[184]);
  assign t[165] = ~(t[78] | t[185]);
  assign t[166] = ~(t[186] & t[105]);
  assign t[167] = ~(t[118] | t[187]);
  assign t[168] = t[163] | t[188];
  assign t[169] = ~(t[233]);
  assign t[16] = ~(t[197] & t[198]);
  assign t[170] = ~(t[226] | t[227]);
  assign t[171] = ~(t[78] | t[189]);
  assign t[172] = ~(t[190] | t[167]);
  assign t[173] = t[195] ? t[159] : t[158];
  assign t[174] = ~(t[234]);
  assign t[175] = ~(t[231] | t[232]);
  assign t[176] = ~(t[136]);
  assign t[177] = ~(t[155] & t[82]);
  assign t[178] = ~(x[4] & t[50]);
  assign t[179] = ~(t[181] & t[82]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[196] | t[198]);
  assign t[181] = ~(x[4] | t[191]);
  assign t[182] = t[195] ? t[119] : t[120];
  assign t[183] = t[195] ? t[192] : t[177];
  assign t[184] = t[195] ? t[158] : t[159];
  assign t[185] = t[195] ? t[177] : t[192];
  assign t[186] = ~(t[48] | t[164]);
  assign t[187] = t[195] ? t[179] : t[158];
  assign t[188] = ~(t[124]);
  assign t[189] = t[195] ? t[178] : t[179];
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[118] | t[193]);
  assign t[191] = ~(t[196]);
  assign t[192] = ~(t[154] & t[198]);
  assign t[193] = t[195] ? t[177] : t[119];
  assign t[194] = t[235] ^ x[2];
  assign t[195] = t[236] ^ x[10];
  assign t[196] = t[237] ^ x[13];
  assign t[197] = t[238] ^ x[16];
  assign t[198] = t[239] ^ x[19];
  assign t[199] = t[240] ^ x[22];
  assign t[19] = t[29] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[241] ^ x[25];
  assign t[201] = t[242] ^ x[27];
  assign t[202] = t[243] ^ x[29];
  assign t[203] = t[244] ^ x[34];
  assign t[204] = t[245] ^ x[37];
  assign t[205] = t[246] ^ x[39];
  assign t[206] = t[247] ^ x[41];
  assign t[207] = t[248] ^ x[44];
  assign t[208] = t[249] ^ x[49];
  assign t[209] = t[250] ^ x[52];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[251] ^ x[54];
  assign t[211] = t[252] ^ x[56];
  assign t[212] = t[253] ^ x[58];
  assign t[213] = t[254] ^ x[62];
  assign t[214] = t[255] ^ x[64];
  assign t[215] = t[256] ^ x[67];
  assign t[216] = t[257] ^ x[71];
  assign t[217] = t[258] ^ x[73];
  assign t[218] = t[259] ^ x[75];
  assign t[219] = t[260] ^ x[77];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[261] ^ x[79];
  assign t[221] = t[262] ^ x[83];
  assign t[222] = t[263] ^ x[85];
  assign t[223] = t[264] ^ x[88];
  assign t[224] = t[265] ^ x[92];
  assign t[225] = t[266] ^ x[94];
  assign t[226] = t[267] ^ x[96];
  assign t[227] = t[268] ^ x[98];
  assign t[228] = t[269] ^ x[100];
  assign t[229] = t[270] ^ x[102];
  assign t[22] = ~(t[21] ^ t[34]);
  assign t[230] = t[271] ^ x[104];
  assign t[231] = t[272] ^ x[106];
  assign t[232] = t[273] ^ x[108];
  assign t[233] = t[274] ^ x[110];
  assign t[234] = t[275] ^ x[112];
  assign t[235] = (x[0] & x[1]);
  assign t[236] = (x[8] & x[9]);
  assign t[237] = (x[11] & x[12]);
  assign t[238] = (x[14] & x[15]);
  assign t[239] = (x[17] & x[18]);
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[240] = (x[20] & x[21]);
  assign t[241] = (x[23] & x[24]);
  assign t[242] = (x[20] & x[26]);
  assign t[243] = (x[20] & x[28]);
  assign t[244] = (x[32] & x[33]);
  assign t[245] = (x[35] & x[36]);
  assign t[246] = (x[23] & x[38]);
  assign t[247] = (x[23] & x[40]);
  assign t[248] = (x[42] & x[43]);
  assign t[249] = (x[47] & x[48]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[50] & x[51]);
  assign t[251] = (x[20] & x[53]);
  assign t[252] = (x[32] & x[55]);
  assign t[253] = (x[32] & x[57]);
  assign t[254] = (x[35] & x[61]);
  assign t[255] = (x[35] & x[63]);
  assign t[256] = (x[65] & x[66]);
  assign t[257] = (x[23] & x[70]);
  assign t[258] = (x[42] & x[72]);
  assign t[259] = (x[42] & x[74]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[260] = (x[47] & x[76]);
  assign t[261] = (x[47] & x[78]);
  assign t[262] = (x[50] & x[82]);
  assign t[263] = (x[50] & x[84]);
  assign t[264] = (x[86] & x[87]);
  assign t[265] = (x[32] & x[91]);
  assign t[266] = (x[35] & x[93]);
  assign t[267] = (x[65] & x[95]);
  assign t[268] = (x[65] & x[97]);
  assign t[269] = (x[42] & x[99]);
  assign t[26] = ~(t[41] ^ t[42]);
  assign t[270] = (x[47] & x[101]);
  assign t[271] = (x[50] & x[103]);
  assign t[272] = (x[86] & x[105]);
  assign t[273] = (x[86] & x[107]);
  assign t[274] = (x[65] & x[109]);
  assign t[275] = (x[86] & x[111]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[29] = ~(t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] & t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[199] | t[54]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[36] = ~(t[43] ^ t[59]);
  assign t[37] = ~(t[60] | t[61]);
  assign t[38] = ~(t[62] ^ t[63]);
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[200] | t[66]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[42] = ~(t[69] ^ t[70]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[44] = ~(t[45] ^ t[73]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[47] = ~(t[197]);
  assign t[48] = ~(t[78] | t[79]);
  assign t[49] = ~(t[80] & t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[196] | t[82]);
  assign t[51] = t[78] & t[195];
  assign t[52] = ~(t[201]);
  assign t[53] = ~(t[202]);
  assign t[54] = ~(t[83] | t[84]);
  assign t[55] = t[197] ? x[31] : x[30];
  assign t[56] = t[85] | t[86];
  assign t[57] = ~(t[87] | t[88]);
  assign t[58] = ~(t[203] | t[89]);
  assign t[59] = ~(t[90] ^ t[91]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[92] | t[93]);
  assign t[61] = ~(t[204] | t[94]);
  assign t[62] = ~(t[95] | t[96]);
  assign t[63] = ~(t[97] ^ t[98]);
  assign t[64] = ~(t[205]);
  assign t[65] = ~(t[206]);
  assign t[66] = ~(t[99] | t[100]);
  assign t[67] = ~(t[101] | t[102]);
  assign t[68] = ~(t[207] | t[103]);
  assign t[69] = t[29] ? x[46] : x[45];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[104] & t[105]);
  assign t[71] = ~(t[106] | t[107]);
  assign t[72] = ~(t[208] | t[108]);
  assign t[73] = ~(t[109] ^ t[110]);
  assign t[74] = ~(t[111] | t[112]);
  assign t[75] = ~(t[209] | t[113]);
  assign t[76] = ~(t[114] | t[115]);
  assign t[77] = ~(t[116] ^ t[117]);
  assign t[78] = ~(t[118]);
  assign t[79] = t[195] ? t[120] : t[119];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121] | t[122]);
  assign t[81] = ~(t[118] & t[123]);
  assign t[82] = ~(t[198]);
  assign t[83] = ~(t[210]);
  assign t[84] = ~(t[201] | t[202]);
  assign t[85] = ~(t[124] & t[31]);
  assign t[86] = ~(t[125] & t[126]);
  assign t[87] = ~(t[211]);
  assign t[88] = ~(t[212]);
  assign t[89] = ~(t[127] | t[128]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[197] ? x[60] : x[59];
  assign t[91] = ~(t[129] & t[130]);
  assign t[92] = ~(t[213]);
  assign t[93] = ~(t[214]);
  assign t[94] = ~(t[131] | t[132]);
  assign t[95] = ~(t[133] | t[134]);
  assign t[96] = ~(t[215] | t[135]);
  assign t[97] = t[197] ? x[69] : x[68];
  assign t[98] = ~(t[129] & t[136]);
  assign t[99] = ~(t[216]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[194];
endmodule

module R1ind162(x, y);
 input [121:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[107] | t[100]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[108] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[31];
  assign t[117] = t[162] ^ x[33];
  assign t[118] = t[163] ^ x[36];
  assign t[119] = t[164] ^ x[39];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[165] ^ x[44];
  assign t[121] = t[166] ^ x[48];
  assign t[122] = t[167] ^ x[50];
  assign t[123] = t[168] ^ x[53];
  assign t[124] = t[169] ^ x[56];
  assign t[125] = t[170] ^ x[61];
  assign t[126] = t[171] ^ x[65];
  assign t[127] = t[172] ^ x[67];
  assign t[128] = t[173] ^ x[69];
  assign t[129] = t[174] ^ x[71];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[73];
  assign t[131] = t[176] ^ x[75];
  assign t[132] = t[177] ^ x[77];
  assign t[133] = t[178] ^ x[79];
  assign t[134] = t[179] ^ x[81];
  assign t[135] = t[180] ^ x[83];
  assign t[136] = t[181] ^ x[85];
  assign t[137] = t[182] ^ x[87];
  assign t[138] = t[183] ^ x[90];
  assign t[139] = t[184] ^ x[92];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[94];
  assign t[141] = t[186] ^ x[97];
  assign t[142] = t[187] ^ x[99];
  assign t[143] = t[188] ^ x[101];
  assign t[144] = t[189] ^ x[103];
  assign t[145] = t[190] ^ x[105];
  assign t[146] = t[191] ^ x[107];
  assign t[147] = t[192] ^ x[109];
  assign t[148] = t[193] ^ x[111];
  assign t[149] = t[194] ^ x[113];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[115];
  assign t[151] = t[196] ^ x[117];
  assign t[152] = t[197] ^ x[119];
  assign t[153] = t[198] ^ x[121];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[20] & x[30]);
  assign t[162] = (x[20] & x[32]);
  assign t[163] = (x[34] & x[35]);
  assign t[164] = (x[37] & x[38]);
  assign t[165] = (x[42] & x[43]);
  assign t[166] = (x[25] & x[47]);
  assign t[167] = (x[25] & x[49]);
  assign t[168] = (x[51] & x[52]);
  assign t[169] = (x[54] & x[55]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[59] & x[60]);
  assign t[171] = (x[20] & x[64]);
  assign t[172] = (x[34] & x[66]);
  assign t[173] = (x[34] & x[68]);
  assign t[174] = (x[37] & x[70]);
  assign t[175] = (x[37] & x[72]);
  assign t[176] = (x[42] & x[74]);
  assign t[177] = (x[42] & x[76]);
  assign t[178] = (x[25] & x[78]);
  assign t[179] = (x[51] & x[80]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[51] & x[82]);
  assign t[181] = (x[54] & x[84]);
  assign t[182] = (x[54] & x[86]);
  assign t[183] = (x[88] & x[89]);
  assign t[184] = (x[59] & x[91]);
  assign t[185] = (x[59] & x[93]);
  assign t[186] = (x[95] & x[96]);
  assign t[187] = (x[34] & x[98]);
  assign t[188] = (x[37] & x[100]);
  assign t[189] = (x[42] & x[102]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[51] & x[104]);
  assign t[191] = (x[54] & x[106]);
  assign t[192] = (x[88] & x[108]);
  assign t[193] = (x[88] & x[110]);
  assign t[194] = (x[59] & x[112]);
  assign t[195] = (x[95] & x[114]);
  assign t[196] = (x[95] & x[116]);
  assign t[197] = (x[88] & x[118]);
  assign t[198] = (x[95] & x[120]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[48] ? x[24] : x[23];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[43];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = t[56] ^ t[35];
  assign t[37] = ~(t[57] & t[58]);
  assign t[38] = t[59] | t[115];
  assign t[39] = t[17] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[69];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[70] | t[45]);
  assign t[48] = ~(t[24]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[73] | t[118];
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = t[76] | t[119];
  assign t[53] = t[112] ? x[41] : x[40];
  assign t[54] = ~(t[77] & t[78]);
  assign t[55] = t[79] | t[120];
  assign t[56] = t[112] ? x[46] : x[45];
  assign t[57] = ~(t[121]);
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[80] | t[57]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[123];
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[124];
  assign t[64] = t[17] ? x[58] : x[57];
  assign t[65] = ~(t[87] & t[88]);
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = t[91] | t[125];
  assign t[68] = t[92] ? x[63] : x[62];
  assign t[69] = ~(t[93] & t[94]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[95] | t[71]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[96] | t[74]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[97] | t[77]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[98] | t[81]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[99] | t[84]);
  assign t[87] = ~(t[100] & t[101]);
  assign t[88] = t[102] | t[138];
  assign t[89] = ~(t[139]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[140]);
  assign t[91] = ~(t[103] | t[89]);
  assign t[92] = ~(t[24]);
  assign t[93] = ~(t[104] & t[105]);
  assign t[94] = t[106] | t[141];
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind163(x, y);
 input [121:0] x;
 output y;

 wire [207:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[144] & t[143]);
  assign t[103] = ~(t[154]);
  assign t[104] = ~(t[146] & t[145]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[114] & t[115]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[116] & t[117]);
  assign t[114] = ~(t[157] & t[156]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[160] & t[159]);
  assign t[117] = ~(t[162]);
  assign t[118] = t[163] ^ x[2];
  assign t[119] = t[164] ^ x[10];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[165] ^ x[13];
  assign t[121] = t[166] ^ x[16];
  assign t[122] = t[167] ^ x[19];
  assign t[123] = t[168] ^ x[22];
  assign t[124] = t[169] ^ x[27];
  assign t[125] = t[170] ^ x[31];
  assign t[126] = t[171] ^ x[33];
  assign t[127] = t[172] ^ x[36];
  assign t[128] = t[173] ^ x[39];
  assign t[129] = t[174] ^ x[44];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[48];
  assign t[131] = t[176] ^ x[50];
  assign t[132] = t[177] ^ x[53];
  assign t[133] = t[178] ^ x[56];
  assign t[134] = t[179] ^ x[61];
  assign t[135] = t[180] ^ x[65];
  assign t[136] = t[181] ^ x[67];
  assign t[137] = t[182] ^ x[69];
  assign t[138] = t[183] ^ x[71];
  assign t[139] = t[184] ^ x[73];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[75];
  assign t[141] = t[186] ^ x[77];
  assign t[142] = t[187] ^ x[79];
  assign t[143] = t[188] ^ x[81];
  assign t[144] = t[189] ^ x[83];
  assign t[145] = t[190] ^ x[85];
  assign t[146] = t[191] ^ x[87];
  assign t[147] = t[192] ^ x[90];
  assign t[148] = t[193] ^ x[92];
  assign t[149] = t[194] ^ x[94];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[97];
  assign t[151] = t[196] ^ x[99];
  assign t[152] = t[197] ^ x[101];
  assign t[153] = t[198] ^ x[103];
  assign t[154] = t[199] ^ x[105];
  assign t[155] = t[200] ^ x[107];
  assign t[156] = t[201] ^ x[109];
  assign t[157] = t[202] ^ x[111];
  assign t[158] = t[203] ^ x[113];
  assign t[159] = t[204] ^ x[115];
  assign t[15] = ~(t[119] & t[120]);
  assign t[160] = t[205] ^ x[117];
  assign t[161] = t[206] ^ x[119];
  assign t[162] = t[207] ^ x[121];
  assign t[163] = (x[0] & x[1]);
  assign t[164] = (x[8] & x[9]);
  assign t[165] = (x[11] & x[12]);
  assign t[166] = (x[14] & x[15]);
  assign t[167] = (x[17] & x[18]);
  assign t[168] = (x[20] & x[21]);
  assign t[169] = (x[25] & x[26]);
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = (x[20] & x[30]);
  assign t[171] = (x[20] & x[32]);
  assign t[172] = (x[34] & x[35]);
  assign t[173] = (x[37] & x[38]);
  assign t[174] = (x[42] & x[43]);
  assign t[175] = (x[25] & x[47]);
  assign t[176] = (x[25] & x[49]);
  assign t[177] = (x[51] & x[52]);
  assign t[178] = (x[54] & x[55]);
  assign t[179] = (x[59] & x[60]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[20] & x[64]);
  assign t[181] = (x[34] & x[66]);
  assign t[182] = (x[34] & x[68]);
  assign t[183] = (x[37] & x[70]);
  assign t[184] = (x[37] & x[72]);
  assign t[185] = (x[42] & x[74]);
  assign t[186] = (x[42] & x[76]);
  assign t[187] = (x[25] & x[78]);
  assign t[188] = (x[51] & x[80]);
  assign t[189] = (x[51] & x[82]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[54] & x[84]);
  assign t[191] = (x[54] & x[86]);
  assign t[192] = (x[88] & x[89]);
  assign t[193] = (x[59] & x[91]);
  assign t[194] = (x[59] & x[93]);
  assign t[195] = (x[95] & x[96]);
  assign t[196] = (x[34] & x[98]);
  assign t[197] = (x[37] & x[100]);
  assign t[198] = (x[42] & x[102]);
  assign t[199] = (x[51] & x[104]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[54] & x[106]);
  assign t[201] = (x[88] & x[108]);
  assign t[202] = (x[88] & x[110]);
  assign t[203] = (x[59] & x[112]);
  assign t[204] = (x[95] & x[114]);
  assign t[205] = (x[95] & x[116]);
  assign t[206] = (x[88] & x[118]);
  assign t[207] = (x[95] & x[120]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[121]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] & t[123]);
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[43];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[35];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = ~(t[58] & t[124]);
  assign t[39] = t[121] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[68];
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[73] & t[127]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = ~(t[76] & t[128]);
  assign t[52] = t[121] ? x[41] : x[40];
  assign t[53] = ~(t[77] & t[78]);
  assign t[54] = ~(t[79] & t[129]);
  assign t[55] = t[121] ? x[46] : x[45];
  assign t[56] = ~(t[130]);
  assign t[57] = ~(t[131]);
  assign t[58] = ~(t[80] & t[81]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[84] & t[132]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[87] & t[133]);
  assign t[63] = t[17] ? x[58] : x[57];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = ~(t[92] & t[134]);
  assign t[67] = t[93] ? x[63] : x[62];
  assign t[68] = ~(t[94] & t[95]);
  assign t[69] = ~(t[126] & t[125]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[135]);
  assign t[71] = ~(t[136]);
  assign t[72] = ~(t[137]);
  assign t[73] = ~(t[96] & t[97]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[139]);
  assign t[76] = ~(t[98] & t[99]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[131] & t[130]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[102] & t[103]);
  assign t[85] = ~(t[145]);
  assign t[86] = ~(t[146]);
  assign t[87] = ~(t[104] & t[105]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[108] & t[147]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[149]);
  assign t[92] = ~(t[109] & t[110]);
  assign t[93] = ~(t[24]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[113] & t[150]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[118];
endmodule

module R1ind164(x, y);
 input [101:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[135] ^ x[10];
  assign t[101] = t[136] ^ x[13];
  assign t[102] = t[137] ^ x[16];
  assign t[103] = t[138] ^ x[19];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[24];
  assign t[106] = t[141] ^ x[29];
  assign t[107] = t[142] ^ x[31];
  assign t[108] = t[143] ^ x[35];
  assign t[109] = t[144] ^ x[38];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] ^ x[40];
  assign t[111] = t[146] ^ x[43];
  assign t[112] = t[147] ^ x[45];
  assign t[113] = t[148] ^ x[50];
  assign t[114] = t[149] ^ x[52];
  assign t[115] = t[150] ^ x[56];
  assign t[116] = t[151] ^ x[59];
  assign t[117] = t[152] ^ x[61];
  assign t[118] = t[153] ^ x[64];
  assign t[119] = t[154] ^ x[66];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[155] ^ x[71];
  assign t[121] = t[156] ^ x[73];
  assign t[122] = t[157] ^ x[77];
  assign t[123] = t[158] ^ x[79];
  assign t[124] = t[159] ^ x[81];
  assign t[125] = t[160] ^ x[83];
  assign t[126] = t[161] ^ x[85];
  assign t[127] = t[162] ^ x[88];
  assign t[128] = t[163] ^ x[90];
  assign t[129] = t[164] ^ x[92];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[165] ^ x[95];
  assign t[131] = t[166] ^ x[97];
  assign t[132] = t[167] ^ x[99];
  assign t[133] = t[168] ^ x[101];
  assign t[134] = (x[0] & x[1]);
  assign t[135] = (x[8] & x[9]);
  assign t[136] = (x[11] & x[12]);
  assign t[137] = (x[14] & x[15]);
  assign t[138] = (x[17] & x[18]);
  assign t[139] = (x[20] & x[21]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[20] & x[23]);
  assign t[141] = (x[27] & x[28]);
  assign t[142] = (x[27] & x[30]);
  assign t[143] = (x[20] & x[34]);
  assign t[144] = (x[36] & x[37]);
  assign t[145] = (x[36] & x[39]);
  assign t[146] = (x[41] & x[42]);
  assign t[147] = (x[41] & x[44]);
  assign t[148] = (x[48] & x[49]);
  assign t[149] = (x[48] & x[51]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[27] & x[55]);
  assign t[151] = (x[57] & x[58]);
  assign t[152] = (x[57] & x[60]);
  assign t[153] = (x[62] & x[63]);
  assign t[154] = (x[62] & x[65]);
  assign t[155] = (x[69] & x[70]);
  assign t[156] = (x[69] & x[72]);
  assign t[157] = (x[36] & x[76]);
  assign t[158] = (x[41] & x[78]);
  assign t[159] = (x[48] & x[80]);
  assign t[15] = ~(t[100] & t[101]);
  assign t[160] = (x[57] & x[82]);
  assign t[161] = (x[62] & x[84]);
  assign t[162] = (x[86] & x[87]);
  assign t[163] = (x[86] & x[89]);
  assign t[164] = (x[69] & x[91]);
  assign t[165] = (x[93] & x[94]);
  assign t[166] = (x[93] & x[96]);
  assign t[167] = (x[86] & x[98]);
  assign t[168] = (x[93] & x[100]);
  assign t[16] = ~(t[102] & t[103]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = t[47] ? x[26] : x[25];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[33];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[43];
  assign t[37] = ~(t[106] & t[56]);
  assign t[38] = ~(t[107] & t[57]);
  assign t[39] = t[58] ? x[33] : x[32];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[68];
  assign t[45] = ~(t[108]);
  assign t[46] = ~(t[108] & t[69]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[109] & t[70]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = t[102] ? x[47] : x[46];
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = ~(t[114] & t[75]);
  assign t[55] = t[102] ? x[54] : x[53];
  assign t[56] = ~(t[115]);
  assign t[57] = ~(t[115] & t[76]);
  assign t[58] = ~(t[24]);
  assign t[59] = ~(t[116] & t[77]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[117] & t[78]);
  assign t[61] = ~(t[118] & t[79]);
  assign t[62] = ~(t[119] & t[80]);
  assign t[63] = t[47] ? x[68] : x[67];
  assign t[64] = ~(t[81] & t[82]);
  assign t[65] = ~(t[120] & t[83]);
  assign t[66] = ~(t[121] & t[84]);
  assign t[67] = t[17] ? x[75] : x[74];
  assign t[68] = ~(t[85] & t[86]);
  assign t[69] = ~(t[104]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[123]);
  assign t[73] = ~(t[123] & t[88]);
  assign t[74] = ~(t[124]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[106]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[125] & t[90]);
  assign t[79] = ~(t[126]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[113]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[116]);
  assign t[91] = ~(t[118]);
  assign t[92] = ~(t[132]);
  assign t[93] = ~(t[132] & t[97]);
  assign t[94] = ~(t[120]);
  assign t[95] = ~(t[133]);
  assign t[96] = ~(t[133] & t[98]);
  assign t[97] = ~(t[127]);
  assign t[98] = ~(t[130]);
  assign t[99] = t[134] ^ x[2];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind165(x, y);
 input [121:0] x;
 output y;

 wire [300:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[233]);
  assign t[101] = ~(t[234]);
  assign t[102] = ~(t[148] | t[149]);
  assign t[103] = t[214] ? x[73] : x[72];
  assign t[104] = t[150] | t[151];
  assign t[105] = ~(t[235]);
  assign t[106] = ~(t[223] | t[224]);
  assign t[107] = ~(t[236]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[152] | t[153]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[139] | t[154]);
  assign t[111] = ~(t[155] | t[84]);
  assign t[112] = ~(t[238]);
  assign t[113] = ~(t[239]);
  assign t[114] = ~(t[156] | t[157]);
  assign t[115] = ~(t[158] | t[159]);
  assign t[116] = ~(t[240] | t[160]);
  assign t[117] = t[29] ? x[88] : x[87];
  assign t[118] = ~(t[161] & t[162]);
  assign t[119] = ~(t[241]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[242]);
  assign t[121] = ~(t[163] | t[164]);
  assign t[122] = ~(t[165] | t[166]);
  assign t[123] = ~(t[243] | t[167]);
  assign t[124] = t[29] ? x[97] : x[96];
  assign t[125] = ~(t[168] & t[169]);
  assign t[126] = ~(t[214]);
  assign t[127] = ~(t[170] & t[171]);
  assign t[128] = ~(t[172] & t[215]);
  assign t[129] = ~(t[215] & t[173]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(x[4] & t[174]);
  assign t[131] = ~(t[175] | t[141]);
  assign t[132] = ~(t[176] & t[177]);
  assign t[133] = t[212] ? t[129] : t[130];
  assign t[134] = ~(t[178]);
  assign t[135] = ~(t[81] | t[179]);
  assign t[136] = t[212] ? t[130] : t[180];
  assign t[137] = ~(t[244]);
  assign t[138] = ~(t[229] | t[230]);
  assign t[139] = ~(t[81] | t[181]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[30] & t[182]);
  assign t[141] = ~(t[126] | t[183]);
  assign t[142] = t[154] | t[134];
  assign t[143] = ~(t[245]);
  assign t[144] = ~(t[231] | t[232]);
  assign t[145] = ~(t[48]);
  assign t[146] = ~(t[150] | t[184]);
  assign t[147] = ~(t[139]);
  assign t[148] = ~(t[246]);
  assign t[149] = ~(t[233] | t[234]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[178] & t[132]);
  assign t[151] = ~(t[110] & t[185]);
  assign t[152] = ~(t[247]);
  assign t[153] = ~(t[236] | t[237]);
  assign t[154] = ~(t[81] | t[186]);
  assign t[155] = ~(t[126] | t[187]);
  assign t[156] = ~(t[248]);
  assign t[157] = ~(t[238] | t[239]);
  assign t[158] = ~(t[249]);
  assign t[159] = ~(t[250]);
  assign t[15] = ~(t[212] & t[213]);
  assign t[160] = ~(t[188] | t[189]);
  assign t[161] = ~(t[155] | t[190]);
  assign t[162] = ~(t[154] | t[191]);
  assign t[163] = ~(t[251]);
  assign t[164] = ~(t[241] | t[242]);
  assign t[165] = ~(t[252]);
  assign t[166] = ~(t[253]);
  assign t[167] = ~(t[192] | t[193]);
  assign t[168] = ~(t[194] | t[195]);
  assign t[169] = ~(t[49] | t[196]);
  assign t[16] = ~(t[214] & t[215]);
  assign t[170] = ~(x[4] | t[213]);
  assign t[171] = ~(t[215]);
  assign t[172] = x[4] & t[213];
  assign t[173] = ~(x[4] | t[197]);
  assign t[174] = ~(t[213] | t[215]);
  assign t[175] = ~(t[126] | t[198]);
  assign t[176] = ~(t[213] | t[171]);
  assign t[177] = t[81] & t[212];
  assign t[178] = ~(t[199] & t[200]);
  assign t[179] = t[212] ? t[201] : t[180];
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[173] & t[171]);
  assign t[181] = t[212] ? t[127] : t[128];
  assign t[182] = ~(t[202] & t[203]);
  assign t[183] = t[212] ? t[180] : t[130];
  assign t[184] = ~(t[204] & t[87]);
  assign t[185] = ~(t[50] | t[196]);
  assign t[186] = t[212] ? t[206] : t[205];
  assign t[187] = t[212] ? t[127] : t[205];
  assign t[188] = ~(t[254]);
  assign t[189] = ~(t[249] | t[250]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[81] | t[207]);
  assign t[191] = ~(t[169] & t[87]);
  assign t[192] = ~(t[255]);
  assign t[193] = ~(t[252] | t[253]);
  assign t[194] = ~(t[161] & t[208]);
  assign t[195] = ~(t[182] & t[87]);
  assign t[196] = ~(t[81] | t[209]);
  assign t[197] = ~(t[213]);
  assign t[198] = t[212] ? t[205] : t[127];
  assign t[199] = ~(t[126] | t[212]);
  assign t[19] = t[29] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = ~(t[129] & t[201]);
  assign t[201] = ~(x[4] & t[176]);
  assign t[202] = t[215] & t[199];
  assign t[203] = t[170] | t[172];
  assign t[204] = ~(t[141]);
  assign t[205] = ~(t[172] & t[171]);
  assign t[206] = ~(t[170] & t[215]);
  assign t[207] = t[212] ? t[180] : t[201];
  assign t[208] = ~(t[126] & t[210]);
  assign t[209] = t[212] ? t[205] : t[206];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = ~(t[130] & t[129]);
  assign t[211] = t[256] ^ x[2];
  assign t[212] = t[257] ^ x[10];
  assign t[213] = t[258] ^ x[13];
  assign t[214] = t[259] ^ x[16];
  assign t[215] = t[260] ^ x[19];
  assign t[216] = t[261] ^ x[22];
  assign t[217] = t[262] ^ x[25];
  assign t[218] = t[263] ^ x[27];
  assign t[219] = t[264] ^ x[29];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[32];
  assign t[221] = t[266] ^ x[37];
  assign t[222] = t[267] ^ x[40];
  assign t[223] = t[268] ^ x[42];
  assign t[224] = t[269] ^ x[44];
  assign t[225] = t[270] ^ x[47];
  assign t[226] = t[271] ^ x[52];
  assign t[227] = t[272] ^ x[55];
  assign t[228] = t[273] ^ x[57];
  assign t[229] = t[274] ^ x[59];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[61];
  assign t[231] = t[276] ^ x[63];
  assign t[232] = t[277] ^ x[65];
  assign t[233] = t[278] ^ x[69];
  assign t[234] = t[279] ^ x[71];
  assign t[235] = t[280] ^ x[75];
  assign t[236] = t[281] ^ x[77];
  assign t[237] = t[282] ^ x[79];
  assign t[238] = t[283] ^ x[81];
  assign t[239] = t[284] ^ x[83];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[86];
  assign t[241] = t[286] ^ x[90];
  assign t[242] = t[287] ^ x[92];
  assign t[243] = t[288] ^ x[95];
  assign t[244] = t[289] ^ x[99];
  assign t[245] = t[290] ^ x[101];
  assign t[246] = t[291] ^ x[103];
  assign t[247] = t[292] ^ x[105];
  assign t[248] = t[293] ^ x[107];
  assign t[249] = t[294] ^ x[109];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = t[295] ^ x[111];
  assign t[251] = t[296] ^ x[113];
  assign t[252] = t[297] ^ x[115];
  assign t[253] = t[298] ^ x[117];
  assign t[254] = t[299] ^ x[119];
  assign t[255] = t[300] ^ x[121];
  assign t[256] = (x[0] & x[1]);
  assign t[257] = (x[8] & x[9]);
  assign t[258] = (x[11] & x[12]);
  assign t[259] = (x[14] & x[15]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[17] & x[18]);
  assign t[261] = (x[20] & x[21]);
  assign t[262] = (x[23] & x[24]);
  assign t[263] = (x[20] & x[26]);
  assign t[264] = (x[20] & x[28]);
  assign t[265] = (x[30] & x[31]);
  assign t[266] = (x[35] & x[36]);
  assign t[267] = (x[38] & x[39]);
  assign t[268] = (x[23] & x[41]);
  assign t[269] = (x[23] & x[43]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[45] & x[46]);
  assign t[271] = (x[50] & x[51]);
  assign t[272] = (x[53] & x[54]);
  assign t[273] = (x[20] & x[56]);
  assign t[274] = (x[30] & x[58]);
  assign t[275] = (x[30] & x[60]);
  assign t[276] = (x[35] & x[62]);
  assign t[277] = (x[35] & x[64]);
  assign t[278] = (x[38] & x[68]);
  assign t[279] = (x[38] & x[70]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[23] & x[74]);
  assign t[281] = (x[45] & x[76]);
  assign t[282] = (x[45] & x[78]);
  assign t[283] = (x[50] & x[80]);
  assign t[284] = (x[50] & x[82]);
  assign t[285] = (x[84] & x[85]);
  assign t[286] = (x[53] & x[89]);
  assign t[287] = (x[53] & x[91]);
  assign t[288] = (x[93] & x[94]);
  assign t[289] = (x[30] & x[98]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[290] = (x[35] & x[100]);
  assign t[291] = (x[38] & x[102]);
  assign t[292] = (x[45] & x[104]);
  assign t[293] = (x[50] & x[106]);
  assign t[294] = (x[84] & x[108]);
  assign t[295] = (x[84] & x[110]);
  assign t[296] = (x[53] & x[112]);
  assign t[297] = (x[93] & x[114]);
  assign t[298] = (x[93] & x[116]);
  assign t[299] = (x[84] & x[118]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[300] = (x[93] & x[120]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51] | t[52]);
  assign t[32] = ~(t[53] | t[54]);
  assign t[33] = ~(t[216] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[58] ^ t[59]);
  assign t[36] = ~(t[60] | t[61]);
  assign t[37] = ~(t[44] ^ t[62]);
  assign t[38] = ~(t[63] | t[64]);
  assign t[39] = ~(t[38] ^ t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[66] | t[67]);
  assign t[41] = ~(t[217] | t[68]);
  assign t[42] = ~(t[69] | t[70]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[45] = ~(t[75] ^ t[76]);
  assign t[46] = ~(t[77] | t[78]);
  assign t[47] = ~(t[79] ^ t[80]);
  assign t[48] = ~(t[214]);
  assign t[49] = ~(t[81] | t[82]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[81] | t[83]);
  assign t[51] = t[84] | t[85];
  assign t[52] = ~(t[86] & t[87]);
  assign t[53] = ~(t[218]);
  assign t[54] = ~(t[219]);
  assign t[55] = ~(t[88] | t[89]);
  assign t[56] = ~(t[90] | t[91]);
  assign t[57] = ~(t[220] | t[92]);
  assign t[58] = t[214] ? x[34] : x[33];
  assign t[59] = ~(t[93] & t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[221] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[100] | t[101]);
  assign t[64] = ~(t[222] | t[102]);
  assign t[65] = ~(t[103] ^ t[104]);
  assign t[66] = ~(t[223]);
  assign t[67] = ~(t[224]);
  assign t[68] = ~(t[105] | t[106]);
  assign t[69] = ~(t[107] | t[108]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[225] | t[109]);
  assign t[71] = t[29] ? x[49] : x[48];
  assign t[72] = ~(t[110] & t[111]);
  assign t[73] = ~(t[112] | t[113]);
  assign t[74] = ~(t[226] | t[114]);
  assign t[75] = ~(t[115] | t[116]);
  assign t[76] = ~(t[117] ^ t[118]);
  assign t[77] = ~(t[119] | t[120]);
  assign t[78] = ~(t[227] | t[121]);
  assign t[79] = ~(t[122] | t[123]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[124] ^ t[125]);
  assign t[81] = ~(t[126]);
  assign t[82] = t[212] ? t[128] : t[127];
  assign t[83] = t[212] ? t[130] : t[129];
  assign t[84] = ~(t[131] & t[132]);
  assign t[85] = ~(t[81] | t[133]);
  assign t[86] = ~(t[134] | t[135]);
  assign t[87] = t[126] | t[136];
  assign t[88] = ~(t[228]);
  assign t[89] = ~(t[218] | t[219]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[229]);
  assign t[91] = ~(t[230]);
  assign t[92] = ~(t[137] | t[138]);
  assign t[93] = ~(t[139] | t[140]);
  assign t[94] = ~(t[141] | t[142]);
  assign t[95] = ~(t[231]);
  assign t[96] = ~(t[232]);
  assign t[97] = ~(t[143] | t[144]);
  assign t[98] = t[145] ? x[67] : x[66];
  assign t[99] = ~(t[146] & t[147]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[211];
endmodule

module R1ind166(x, y);
 input [85:0] x;
 output y;

 wire [142:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[65];
  assign t[101] = t[133] ^ x[67];
  assign t[102] = t[134] ^ x[69];
  assign t[103] = t[135] ^ x[71];
  assign t[104] = t[136] ^ x[73];
  assign t[105] = t[137] ^ x[75];
  assign t[106] = t[138] ^ x[77];
  assign t[107] = t[139] ^ x[79];
  assign t[108] = t[140] ^ x[81];
  assign t[109] = t[141] ^ x[83];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[85];
  assign t[111] = (x[0] & x[1]);
  assign t[112] = (x[8] & x[9]);
  assign t[113] = (x[11] & x[12]);
  assign t[114] = (x[14] & x[15]);
  assign t[115] = (x[17] & x[18]);
  assign t[116] = (x[20] & x[21]);
  assign t[117] = (x[0] & x[23]);
  assign t[118] = (x[20] & x[27]);
  assign t[119] = (x[20] & x[29]);
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = (x[31] & x[32]);
  assign t[121] = (x[36] & x[37]);
  assign t[122] = (x[0] & x[41]);
  assign t[123] = (x[43] & x[44]);
  assign t[124] = (x[20] & x[46]);
  assign t[125] = (x[31] & x[48]);
  assign t[126] = (x[31] & x[50]);
  assign t[127] = (x[52] & x[53]);
  assign t[128] = (x[36] & x[55]);
  assign t[129] = (x[36] & x[57]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[130] = (x[59] & x[60]);
  assign t[131] = (x[0] & x[62]);
  assign t[132] = (x[43] & x[64]);
  assign t[133] = (x[43] & x[66]);
  assign t[134] = (x[31] & x[68]);
  assign t[135] = (x[52] & x[70]);
  assign t[136] = (x[52] & x[72]);
  assign t[137] = (x[36] & x[74]);
  assign t[138] = (x[59] & x[76]);
  assign t[139] = (x[59] & x[78]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = (x[43] & x[80]);
  assign t[141] = (x[52] & x[82]);
  assign t[142] = (x[59] & x[84]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[80] & t[81]);
  assign t[16] = ~(t[82] & t[83]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[82]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[36] & t[37]);
  assign t[27] = t[38] | t[84];
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = t[41] ^ t[42];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[43] & t[44]);
  assign t[31] = t[45] ^ t[46];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] | t[85];
  assign t[34] = t[17] ? x[26] : x[25];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = ~(t[86]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[52] | t[36]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[55] | t[88];
  assign t[41] = t[17] ? x[35] : x[34];
  assign t[42] = ~(t[56] & t[57]);
  assign t[43] = ~(t[58] & t[59]);
  assign t[44] = t[60] | t[89];
  assign t[45] = t[61] ? x[40] : x[39];
  assign t[46] = ~(t[62] & t[63]);
  assign t[47] = ~(t[79]);
  assign t[48] = ~(t[90]);
  assign t[49] = ~(t[64] | t[47]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[65] & t[66]);
  assign t[51] = t[67] | t[91];
  assign t[52] = ~(t[92]);
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[68] | t[53]);
  assign t[56] = ~(t[69] & t[70]);
  assign t[57] = t[71] | t[95];
  assign t[58] = ~(t[96]);
  assign t[59] = ~(t[97]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[72] | t[58]);
  assign t[61] = ~(t[23]);
  assign t[62] = ~(t[73] & t[74]);
  assign t[63] = t[75] | t[98];
  assign t[64] = ~(t[99]);
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[76] | t[65]);
  assign t[68] = ~(t[102]);
  assign t[69] = ~(t[103]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[77] | t[69]);
  assign t[72] = ~(t[105]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[78] | t[73]);
  assign t[76] = ~(t[108]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = t[111] ^ x[2];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[112] ^ x[10];
  assign t[81] = t[113] ^ x[13];
  assign t[82] = t[114] ^ x[16];
  assign t[83] = t[115] ^ x[19];
  assign t[84] = t[116] ^ x[22];
  assign t[85] = t[117] ^ x[24];
  assign t[86] = t[118] ^ x[28];
  assign t[87] = t[119] ^ x[30];
  assign t[88] = t[120] ^ x[33];
  assign t[89] = t[121] ^ x[38];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[122] ^ x[42];
  assign t[91] = t[123] ^ x[45];
  assign t[92] = t[124] ^ x[47];
  assign t[93] = t[125] ^ x[49];
  assign t[94] = t[126] ^ x[51];
  assign t[95] = t[127] ^ x[54];
  assign t[96] = t[128] ^ x[56];
  assign t[97] = t[129] ^ x[58];
  assign t[98] = t[130] ^ x[61];
  assign t[99] = t[131] ^ x[63];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[79];
endmodule

module R1ind167(x, y);
 input [85:0] x;
 output y;

 wire [149:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[49];
  assign t[101] = t[133] ^ x[51];
  assign t[102] = t[134] ^ x[53];
  assign t[103] = t[135] ^ x[56];
  assign t[104] = t[136] ^ x[58];
  assign t[105] = t[137] ^ x[60];
  assign t[106] = t[138] ^ x[63];
  assign t[107] = t[139] ^ x[65];
  assign t[108] = t[140] ^ x[67];
  assign t[109] = t[141] ^ x[69];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[71];
  assign t[111] = t[143] ^ x[73];
  assign t[112] = t[144] ^ x[75];
  assign t[113] = t[145] ^ x[77];
  assign t[114] = t[146] ^ x[79];
  assign t[115] = t[147] ^ x[81];
  assign t[116] = t[148] ^ x[83];
  assign t[117] = t[149] ^ x[85];
  assign t[118] = (x[0] & x[1]);
  assign t[119] = (x[8] & x[9]);
  assign t[11] = t[87] ? x[6] : x[7];
  assign t[120] = (x[11] & x[12]);
  assign t[121] = (x[14] & x[15]);
  assign t[122] = (x[17] & x[18]);
  assign t[123] = (x[20] & x[21]);
  assign t[124] = (x[0] & x[23]);
  assign t[125] = (x[20] & x[27]);
  assign t[126] = (x[20] & x[29]);
  assign t[127] = (x[31] & x[32]);
  assign t[128] = (x[36] & x[37]);
  assign t[129] = (x[0] & x[41]);
  assign t[12] = ~(t[17] ^ t[14]);
  assign t[130] = (x[0] & x[43]);
  assign t[131] = (x[45] & x[46]);
  assign t[132] = (x[20] & x[48]);
  assign t[133] = (x[31] & x[50]);
  assign t[134] = (x[31] & x[52]);
  assign t[135] = (x[54] & x[55]);
  assign t[136] = (x[36] & x[57]);
  assign t[137] = (x[36] & x[59]);
  assign t[138] = (x[61] & x[62]);
  assign t[139] = (x[45] & x[64]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (x[45] & x[66]);
  assign t[141] = (x[31] & x[68]);
  assign t[142] = (x[54] & x[70]);
  assign t[143] = (x[54] & x[72]);
  assign t[144] = (x[36] & x[74]);
  assign t[145] = (x[61] & x[76]);
  assign t[146] = (x[61] & x[78]);
  assign t[147] = (x[45] & x[80]);
  assign t[148] = (x[54] & x[82]);
  assign t[149] = (x[61] & x[84]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[15] = ~(t[88] & t[89]);
  assign t[16] = ~(t[87] & t[90]);
  assign t[17] = x[4] ? t[23] : t[22];
  assign t[18] = ~(t[24] & t[25]);
  assign t[19] = t[11] ^ t[22];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = x[4] ? t[27] : t[26];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = t[32] ^ t[33];
  assign t[24] = ~(t[34] & t[35]);
  assign t[25] = ~(t[36] & t[91]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[27] = t[39] ^ t[40];
  assign t[28] = ~(t[41] & t[42]);
  assign t[29] = t[43] ^ t[44];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[31] = ~(t[47] & t[92]);
  assign t[32] = t[48] ? x[26] : x[25];
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = ~(t[93]);
  assign t[35] = ~(t[94]);
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[53] & t[54]);
  assign t[38] = ~(t[55] & t[95]);
  assign t[39] = t[48] ? x[35] : x[34];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[56] & t[57]);
  assign t[41] = ~(t[58] & t[59]);
  assign t[42] = ~(t[60] & t[96]);
  assign t[43] = t[61] ? x[40] : x[39];
  assign t[44] = ~(t[62] & t[63]);
  assign t[45] = ~(t[97]);
  assign t[46] = ~(t[98]);
  assign t[47] = ~(t[64] & t[65]);
  assign t[48] = ~(t[66]);
  assign t[49] = ~(t[67] & t[68]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[69] & t[99]);
  assign t[51] = ~(t[94] & t[93]);
  assign t[52] = ~(t[100]);
  assign t[53] = ~(t[101]);
  assign t[54] = ~(t[102]);
  assign t[55] = ~(t[70] & t[71]);
  assign t[56] = ~(t[72] & t[73]);
  assign t[57] = ~(t[74] & t[103]);
  assign t[58] = ~(t[104]);
  assign t[59] = ~(t[105]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[75] & t[76]);
  assign t[61] = ~(t[66]);
  assign t[62] = ~(t[77] & t[78]);
  assign t[63] = ~(t[79] & t[106]);
  assign t[64] = ~(t[98] & t[97]);
  assign t[65] = ~(t[86]);
  assign t[66] = ~(t[87]);
  assign t[67] = ~(t[107]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[80] & t[81]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[102] & t[101]);
  assign t[71] = ~(t[109]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[82] & t[83]);
  assign t[75] = ~(t[105] & t[104]);
  assign t[76] = ~(t[112]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[84] & t[85]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[108] & t[107]);
  assign t[81] = ~(t[115]);
  assign t[82] = ~(t[111] & t[110]);
  assign t[83] = ~(t[116]);
  assign t[84] = ~(t[114] & t[113]);
  assign t[85] = ~(t[117]);
  assign t[86] = t[118] ^ x[2];
  assign t[87] = t[119] ^ x[10];
  assign t[88] = t[120] ^ x[13];
  assign t[89] = t[121] ^ x[16];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[122] ^ x[19];
  assign t[91] = t[123] ^ x[22];
  assign t[92] = t[124] ^ x[24];
  assign t[93] = t[125] ^ x[28];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[33];
  assign t[96] = t[128] ^ x[38];
  assign t[97] = t[129] ^ x[42];
  assign t[98] = t[130] ^ x[44];
  assign t[99] = t[131] ^ x[47];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[86];
endmodule

module R1ind168(x, y);
 input [73:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = (x[8] & x[9]);
  assign t[101] = (x[11] & x[12]);
  assign t[102] = (x[14] & x[15]);
  assign t[103] = (x[17] & x[18]);
  assign t[104] = (x[20] & x[21]);
  assign t[105] = (x[20] & x[23]);
  assign t[106] = (x[0] & x[25]);
  assign t[107] = (x[0] & x[27]);
  assign t[108] = (x[20] & x[31]);
  assign t[109] = (x[33] & x[34]);
  assign t[10] = ~(x[3]);
  assign t[110] = (x[33] & x[36]);
  assign t[111] = (x[40] & x[41]);
  assign t[112] = (x[40] & x[43]);
  assign t[113] = (x[0] & x[47]);
  assign t[114] = (x[49] & x[50]);
  assign t[115] = (x[49] & x[52]);
  assign t[116] = (x[33] & x[54]);
  assign t[117] = (x[56] & x[57]);
  assign t[118] = (x[56] & x[59]);
  assign t[119] = (x[40] & x[61]);
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = (x[63] & x[64]);
  assign t[121] = (x[63] & x[66]);
  assign t[122] = (x[49] & x[68]);
  assign t[123] = (x[56] & x[70]);
  assign t[124] = (x[63] & x[72]);
  assign t[12] = ~(t[18] ^ t[14]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[74] & t[75]);
  assign t[16] = ~(t[76] & t[77]);
  assign t[17] = ~(t[23]);
  assign t[18] = x[4] ? t[25] : t[24];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[11] ^ t[24];
  assign t[21] = x[4] ? t[29] : t[28];
  assign t[22] = x[4] ? t[31] : t[30];
  assign t[23] = ~(t[76]);
  assign t[24] = ~(t[32] & t[33]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[78] & t[36]);
  assign t[27] = ~(t[79] & t[37]);
  assign t[28] = ~(t[38] & t[39]);
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[42] & t[43]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[80] & t[46]);
  assign t[33] = ~(t[81] & t[47]);
  assign t[34] = t[48] ? x[30] : x[29];
  assign t[35] = ~(t[49] & t[50]);
  assign t[36] = ~(t[82]);
  assign t[37] = ~(t[82] & t[51]);
  assign t[38] = ~(t[83] & t[52]);
  assign t[39] = ~(t[84] & t[53]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[54] ? x[39] : x[38];
  assign t[41] = ~(t[55] & t[56]);
  assign t[42] = ~(t[85] & t[57]);
  assign t[43] = ~(t[86] & t[58]);
  assign t[44] = t[48] ? x[46] : x[45];
  assign t[45] = ~(t[59] & t[60]);
  assign t[46] = ~(t[87]);
  assign t[47] = ~(t[87] & t[61]);
  assign t[48] = ~(t[23]);
  assign t[49] = ~(t[88] & t[62]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[89] & t[63]);
  assign t[51] = ~(t[78]);
  assign t[52] = ~(t[90]);
  assign t[53] = ~(t[90] & t[64]);
  assign t[54] = ~(t[23]);
  assign t[55] = ~(t[91] & t[65]);
  assign t[56] = ~(t[92] & t[66]);
  assign t[57] = ~(t[93]);
  assign t[58] = ~(t[93] & t[67]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] & t[69]);
  assign t[61] = ~(t[80]);
  assign t[62] = ~(t[96]);
  assign t[63] = ~(t[96] & t[70]);
  assign t[64] = ~(t[83]);
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[97] & t[71]);
  assign t[67] = ~(t[85]);
  assign t[68] = ~(t[98]);
  assign t[69] = ~(t[98] & t[72]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[88]);
  assign t[71] = ~(t[91]);
  assign t[72] = ~(t[94]);
  assign t[73] = t[99] ^ x[2];
  assign t[74] = t[100] ^ x[10];
  assign t[75] = t[101] ^ x[13];
  assign t[76] = t[102] ^ x[16];
  assign t[77] = t[103] ^ x[19];
  assign t[78] = t[104] ^ x[22];
  assign t[79] = t[105] ^ x[24];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[106] ^ x[26];
  assign t[81] = t[107] ^ x[28];
  assign t[82] = t[108] ^ x[32];
  assign t[83] = t[109] ^ x[35];
  assign t[84] = t[110] ^ x[37];
  assign t[85] = t[111] ^ x[42];
  assign t[86] = t[112] ^ x[44];
  assign t[87] = t[113] ^ x[48];
  assign t[88] = t[114] ^ x[51];
  assign t[89] = t[115] ^ x[53];
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[116] ^ x[55];
  assign t[91] = t[117] ^ x[58];
  assign t[92] = t[118] ^ x[60];
  assign t[93] = t[119] ^ x[62];
  assign t[94] = t[120] ^ x[65];
  assign t[95] = t[121] ^ x[67];
  assign t[96] = t[122] ^ x[69];
  assign t[97] = t[123] ^ x[71];
  assign t[98] = t[124] ^ x[73];
  assign t[99] = (x[0] & x[1]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[73];
endmodule

module R1ind169(x, y);
 input [85:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[184]);
  assign t[101] = ~(t[176] | t[177]);
  assign t[102] = ~(t[185]);
  assign t[103] = ~(t[186]);
  assign t[104] = ~(t[125] | t[126]);
  assign t[105] = ~(t[42] | t[127]);
  assign t[106] = ~(t[41] | t[128]);
  assign t[107] = ~(t[187]);
  assign t[108] = ~(t[179] | t[180]);
  assign t[109] = ~(t[188]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[189]);
  assign t[111] = ~(t[129] | t[130]);
  assign t[112] = ~(t[131] | t[132]);
  assign t[113] = ~(t[116] | t[133]);
  assign t[114] = ~(t[190]);
  assign t[115] = ~(t[182] | t[183]);
  assign t[116] = ~(t[62] | t[134]);
  assign t[117] = ~(t[62] | t[135]);
  assign t[118] = t[43] | t[136];
  assign t[119] = ~(t[137] & t[138]);
  assign t[11] = ~(t[17] ^ t[14]);
  assign t[120] = x[4] & t[163];
  assign t[121] = ~(x[4] | t[163]);
  assign t[122] = ~(t[165]);
  assign t[123] = t[162] ? t[94] : t[93];
  assign t[124] = t[162] ? t[140] : t[139];
  assign t[125] = ~(t[191]);
  assign t[126] = ~(t[185] | t[186]);
  assign t[127] = ~(t[62] | t[141]);
  assign t[128] = ~(t[113] & t[138]);
  assign t[129] = ~(t[192]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[188] | t[189]);
  assign t[131] = ~(t[105] & t[142]);
  assign t[132] = ~(t[143] & t[138]);
  assign t[133] = ~(t[62] | t[144]);
  assign t[134] = t[162] ? t[92] : t[93];
  assign t[135] = t[162] ? t[139] : t[145];
  assign t[136] = ~(t[62] | t[146]);
  assign t[137] = ~(t[147] | t[148]);
  assign t[138] = t[65] | t[149];
  assign t[139] = ~(x[4] & t[150]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = ~(t[151] & t[122]);
  assign t[141] = t[162] ? t[140] : t[152];
  assign t[142] = ~(t[65] & t[153]);
  assign t[143] = ~(t[154] & t[155]);
  assign t[144] = t[162] ? t[94] : t[95];
  assign t[145] = ~(t[165] & t[151]);
  assign t[146] = t[162] ? t[145] : t[139];
  assign t[147] = ~(t[156]);
  assign t[148] = ~(t[62] | t[157]);
  assign t[149] = t[162] ? t[139] : t[140];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = ~(t[163] | t[165]);
  assign t[151] = ~(x[4] | t[158]);
  assign t[152] = ~(x[4] & t[98]);
  assign t[153] = ~(t[139] & t[145]);
  assign t[154] = t[165] & t[159];
  assign t[155] = t[121] | t[120];
  assign t[156] = ~(t[159] & t[160]);
  assign t[157] = t[162] ? t[152] : t[140];
  assign t[158] = ~(t[163]);
  assign t[159] = ~(t[65] | t[162]);
  assign t[15] = ~(t[162] & t[163]);
  assign t[160] = ~(t[145] & t[152]);
  assign t[161] = t[193] ^ x[2];
  assign t[162] = t[194] ^ x[10];
  assign t[163] = t[195] ^ x[13];
  assign t[164] = t[196] ^ x[16];
  assign t[165] = t[197] ^ x[19];
  assign t[166] = t[198] ^ x[22];
  assign t[167] = t[199] ^ x[24];
  assign t[168] = t[200] ^ x[26];
  assign t[169] = t[201] ^ x[28];
  assign t[16] = ~(t[164] & t[165]);
  assign t[170] = t[202] ^ x[31];
  assign t[171] = t[203] ^ x[34];
  assign t[172] = t[204] ^ x[36];
  assign t[173] = t[205] ^ x[38];
  assign t[174] = t[206] ^ x[41];
  assign t[175] = t[207] ^ x[45];
  assign t[176] = t[208] ^ x[47];
  assign t[177] = t[209] ^ x[49];
  assign t[178] = t[210] ^ x[52];
  assign t[179] = t[211] ^ x[56];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[180] = t[212] ^ x[58];
  assign t[181] = t[213] ^ x[61];
  assign t[182] = t[214] ^ x[65];
  assign t[183] = t[215] ^ x[67];
  assign t[184] = t[216] ^ x[69];
  assign t[185] = t[217] ^ x[71];
  assign t[186] = t[218] ^ x[73];
  assign t[187] = t[219] ^ x[75];
  assign t[188] = t[220] ^ x[77];
  assign t[189] = t[221] ^ x[79];
  assign t[18] = t[26] ? x[6] : x[7];
  assign t[190] = t[222] ^ x[81];
  assign t[191] = t[223] ^ x[83];
  assign t[192] = t[224] ^ x[85];
  assign t[193] = (x[0] & x[1]);
  assign t[194] = (x[8] & x[9]);
  assign t[195] = (x[11] & x[12]);
  assign t[196] = (x[14] & x[15]);
  assign t[197] = (x[17] & x[18]);
  assign t[198] = (x[20] & x[21]);
  assign t[199] = (x[0] & x[23]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[20] & x[25]);
  assign t[201] = (x[20] & x[27]);
  assign t[202] = (x[29] & x[30]);
  assign t[203] = (x[32] & x[33]);
  assign t[204] = (x[0] & x[35]);
  assign t[205] = (x[0] & x[37]);
  assign t[206] = (x[39] & x[40]);
  assign t[207] = (x[20] & x[44]);
  assign t[208] = (x[29] & x[46]);
  assign t[209] = (x[29] & x[48]);
  assign t[20] = ~(t[29] | t[30]);
  assign t[210] = (x[50] & x[51]);
  assign t[211] = (x[32] & x[55]);
  assign t[212] = (x[32] & x[57]);
  assign t[213] = (x[59] & x[60]);
  assign t[214] = (x[39] & x[64]);
  assign t[215] = (x[39] & x[66]);
  assign t[216] = (x[29] & x[68]);
  assign t[217] = (x[50] & x[70]);
  assign t[218] = (x[50] & x[72]);
  assign t[219] = (x[32] & x[74]);
  assign t[21] = ~(t[24] ^ t[12]);
  assign t[220] = (x[59] & x[76]);
  assign t[221] = (x[59] & x[78]);
  assign t[222] = (x[39] & x[80]);
  assign t[223] = (x[50] & x[82]);
  assign t[224] = (x[59] & x[84]);
  assign t[22] = x[4] ? t[32] : t[31];
  assign t[23] = x[4] ? t[34] : t[33];
  assign t[24] = ~(t[35] | t[36]);
  assign t[25] = ~(t[37] ^ t[38]);
  assign t[26] = ~(t[39]);
  assign t[27] = ~(t[40] | t[41]);
  assign t[28] = ~(t[42] | t[43]);
  assign t[29] = ~(t[44] | t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[166] | t[46]);
  assign t[31] = ~(t[47] | t[48]);
  assign t[32] = ~(t[49] ^ t[50]);
  assign t[33] = ~(t[51] | t[52]);
  assign t[34] = ~(t[53] ^ t[54]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[167] | t[57]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = ~(t[60] ^ t[61]);
  assign t[39] = ~(t[164]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[62] | t[63]);
  assign t[41] = ~(t[62] | t[64]);
  assign t[42] = ~(t[65] | t[66]);
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = ~(t[168]);
  assign t[45] = ~(t[169]);
  assign t[46] = ~(t[69] | t[70]);
  assign t[47] = ~(t[71] | t[72]);
  assign t[48] = ~(t[170] | t[73]);
  assign t[49] = ~(t[74] | t[75]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[76] ^ t[77]);
  assign t[51] = ~(t[78] | t[79]);
  assign t[52] = ~(t[171] | t[80]);
  assign t[53] = ~(t[81] | t[82]);
  assign t[54] = ~(t[83] ^ t[84]);
  assign t[55] = ~(t[172]);
  assign t[56] = ~(t[173]);
  assign t[57] = ~(t[85] | t[86]);
  assign t[58] = ~(t[87] | t[88]);
  assign t[59] = ~(t[174] | t[89]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[26] ? x[43] : x[42];
  assign t[61] = ~(t[90] & t[91]);
  assign t[62] = ~(t[65]);
  assign t[63] = t[162] ? t[93] : t[92];
  assign t[64] = t[162] ? t[95] : t[94];
  assign t[65] = ~(t[164]);
  assign t[66] = t[162] ? t[93] : t[94];
  assign t[67] = ~(t[96] | t[97]);
  assign t[68] = ~(t[98] & t[99]);
  assign t[69] = ~(t[175]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[168] | t[169]);
  assign t[71] = ~(t[176]);
  assign t[72] = ~(t[177]);
  assign t[73] = ~(t[100] | t[101]);
  assign t[74] = ~(t[102] | t[103]);
  assign t[75] = ~(t[178] | t[104]);
  assign t[76] = t[26] ? x[54] : x[53];
  assign t[77] = ~(t[105] & t[106]);
  assign t[78] = ~(t[179]);
  assign t[79] = ~(t[180]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[107] | t[108]);
  assign t[81] = ~(t[109] | t[110]);
  assign t[82] = ~(t[181] | t[111]);
  assign t[83] = t[26] ? x[63] : x[62];
  assign t[84] = ~(t[112] & t[113]);
  assign t[85] = ~(t[161]);
  assign t[86] = ~(t[172] | t[173]);
  assign t[87] = ~(t[182]);
  assign t[88] = ~(t[183]);
  assign t[89] = ~(t[114] | t[115]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[116] | t[117]);
  assign t[91] = ~(t[118] | t[119]);
  assign t[92] = ~(t[120] & t[165]);
  assign t[93] = ~(t[121] & t[122]);
  assign t[94] = ~(t[120] & t[122]);
  assign t[95] = ~(t[121] & t[165]);
  assign t[96] = ~(t[65] | t[123]);
  assign t[97] = ~(t[65] | t[124]);
  assign t[98] = ~(t[163] | t[122]);
  assign t[99] = t[62] & t[162];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[161];
endmodule

module R1ind170(x, y);
 input [112:0] x;
 output y;

 wire [183:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = t[143] ^ x[2];
  assign t[103] = t[144] ^ x[10];
  assign t[104] = t[145] ^ x[13];
  assign t[105] = t[146] ^ x[16];
  assign t[106] = t[147] ^ x[19];
  assign t[107] = t[148] ^ x[22];
  assign t[108] = t[149] ^ x[27];
  assign t[109] = t[150] ^ x[31];
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[33];
  assign t[111] = t[152] ^ x[36];
  assign t[112] = t[153] ^ x[41];
  assign t[113] = t[154] ^ x[45];
  assign t[114] = t[155] ^ x[47];
  assign t[115] = t[156] ^ x[50];
  assign t[116] = t[157] ^ x[53];
  assign t[117] = t[158] ^ x[58];
  assign t[118] = t[159] ^ x[62];
  assign t[119] = t[160] ^ x[64];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[66];
  assign t[121] = t[162] ^ x[68];
  assign t[122] = t[163] ^ x[70];
  assign t[123] = t[164] ^ x[73];
  assign t[124] = t[165] ^ x[75];
  assign t[125] = t[166] ^ x[77];
  assign t[126] = t[167] ^ x[79];
  assign t[127] = t[168] ^ x[81];
  assign t[128] = t[169] ^ x[83];
  assign t[129] = t[170] ^ x[86];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[88];
  assign t[131] = t[172] ^ x[90];
  assign t[132] = t[173] ^ x[92];
  assign t[133] = t[174] ^ x[94];
  assign t[134] = t[175] ^ x[96];
  assign t[135] = t[176] ^ x[98];
  assign t[136] = t[177] ^ x[100];
  assign t[137] = t[178] ^ x[102];
  assign t[138] = t[179] ^ x[104];
  assign t[139] = t[180] ^ x[106];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[108];
  assign t[141] = t[182] ^ x[110];
  assign t[142] = t[183] ^ x[112];
  assign t[143] = (x[0] & x[1]);
  assign t[144] = (x[8] & x[9]);
  assign t[145] = (x[11] & x[12]);
  assign t[146] = (x[14] & x[15]);
  assign t[147] = (x[17] & x[18]);
  assign t[148] = (x[20] & x[21]);
  assign t[149] = (x[25] & x[26]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[20] & x[30]);
  assign t[151] = (x[20] & x[32]);
  assign t[152] = (x[34] & x[35]);
  assign t[153] = (x[39] & x[40]);
  assign t[154] = (x[25] & x[44]);
  assign t[155] = (x[25] & x[46]);
  assign t[156] = (x[48] & x[49]);
  assign t[157] = (x[51] & x[52]);
  assign t[158] = (x[56] & x[57]);
  assign t[159] = (x[20] & x[61]);
  assign t[15] = ~(t[103] & t[104]);
  assign t[160] = (x[34] & x[63]);
  assign t[161] = (x[34] & x[65]);
  assign t[162] = (x[39] & x[67]);
  assign t[163] = (x[39] & x[69]);
  assign t[164] = (x[71] & x[72]);
  assign t[165] = (x[25] & x[74]);
  assign t[166] = (x[48] & x[76]);
  assign t[167] = (x[48] & x[78]);
  assign t[168] = (x[51] & x[80]);
  assign t[169] = (x[51] & x[82]);
  assign t[16] = ~(t[105] & t[106]);
  assign t[170] = (x[84] & x[85]);
  assign t[171] = (x[56] & x[87]);
  assign t[172] = (x[56] & x[89]);
  assign t[173] = (x[34] & x[91]);
  assign t[174] = (x[39] & x[93]);
  assign t[175] = (x[71] & x[95]);
  assign t[176] = (x[71] & x[97]);
  assign t[177] = (x[48] & x[99]);
  assign t[178] = (x[51] & x[101]);
  assign t[179] = (x[84] & x[103]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[84] & x[105]);
  assign t[181] = (x[56] & x[107]);
  assign t[182] = (x[71] & x[109]);
  assign t[183] = (x[84] & x[111]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[105]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] | t[107];
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[42];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[53];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] | t[108];
  assign t[38] = t[57] ? x[29] : x[28];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[63];
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[40];
  assign t[44] = ~(t[109]);
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[67] | t[44]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = t[70] | t[111];
  assign t[49] = t[71] ? x[38] : x[37];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[112];
  assign t[52] = t[17] ? x[43] : x[42];
  assign t[53] = ~(t[75] & t[76]);
  assign t[54] = ~(t[113]);
  assign t[55] = ~(t[114]);
  assign t[56] = ~(t[77] | t[54]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[78] & t[79]);
  assign t[59] = t[80] | t[115];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[116];
  assign t[62] = t[57] ? x[55] : x[54];
  assign t[63] = ~(t[84] & t[85]);
  assign t[64] = ~(t[86] & t[87]);
  assign t[65] = t[88] | t[117];
  assign t[66] = t[57] ? x[60] : x[59];
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[89] | t[68]);
  assign t[71] = ~(t[24]);
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[90] | t[72]);
  assign t[75] = ~(t[91] & t[92]);
  assign t[76] = t[93] | t[123];
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[94] | t[78]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[95] | t[81]);
  assign t[84] = ~(t[96] & t[97]);
  assign t[85] = t[98] | t[129];
  assign t[86] = ~(t[130]);
  assign t[87] = ~(t[131]);
  assign t[88] = ~(t[99] | t[86]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[100] | t[91]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[101] | t[96]);
  assign t[99] = ~(t[140]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[102];
endmodule

module R1ind171(x, y);
 input [112:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[109] & t[110]);
  assign t[105] = ~(t[140] & t[139]);
  assign t[106] = ~(t[149]);
  assign t[107] = ~(t[144] & t[143]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[148] & t[147]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[151]);
  assign t[111] = t[152] ^ x[2];
  assign t[112] = t[153] ^ x[10];
  assign t[113] = t[154] ^ x[13];
  assign t[114] = t[155] ^ x[16];
  assign t[115] = t[156] ^ x[19];
  assign t[116] = t[157] ^ x[22];
  assign t[117] = t[158] ^ x[27];
  assign t[118] = t[159] ^ x[31];
  assign t[119] = t[160] ^ x[33];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[36];
  assign t[121] = t[162] ^ x[41];
  assign t[122] = t[163] ^ x[45];
  assign t[123] = t[164] ^ x[47];
  assign t[124] = t[165] ^ x[50];
  assign t[125] = t[166] ^ x[53];
  assign t[126] = t[167] ^ x[58];
  assign t[127] = t[168] ^ x[62];
  assign t[128] = t[169] ^ x[64];
  assign t[129] = t[170] ^ x[66];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[171] ^ x[68];
  assign t[131] = t[172] ^ x[70];
  assign t[132] = t[173] ^ x[73];
  assign t[133] = t[174] ^ x[75];
  assign t[134] = t[175] ^ x[77];
  assign t[135] = t[176] ^ x[79];
  assign t[136] = t[177] ^ x[81];
  assign t[137] = t[178] ^ x[83];
  assign t[138] = t[179] ^ x[86];
  assign t[139] = t[180] ^ x[88];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[181] ^ x[90];
  assign t[141] = t[182] ^ x[92];
  assign t[142] = t[183] ^ x[94];
  assign t[143] = t[184] ^ x[96];
  assign t[144] = t[185] ^ x[98];
  assign t[145] = t[186] ^ x[100];
  assign t[146] = t[187] ^ x[102];
  assign t[147] = t[188] ^ x[104];
  assign t[148] = t[189] ^ x[106];
  assign t[149] = t[190] ^ x[108];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[191] ^ x[110];
  assign t[151] = t[192] ^ x[112];
  assign t[152] = (x[0] & x[1]);
  assign t[153] = (x[8] & x[9]);
  assign t[154] = (x[11] & x[12]);
  assign t[155] = (x[14] & x[15]);
  assign t[156] = (x[17] & x[18]);
  assign t[157] = (x[20] & x[21]);
  assign t[158] = (x[25] & x[26]);
  assign t[159] = (x[20] & x[30]);
  assign t[15] = ~(t[112] & t[113]);
  assign t[160] = (x[20] & x[32]);
  assign t[161] = (x[34] & x[35]);
  assign t[162] = (x[39] & x[40]);
  assign t[163] = (x[25] & x[44]);
  assign t[164] = (x[25] & x[46]);
  assign t[165] = (x[48] & x[49]);
  assign t[166] = (x[51] & x[52]);
  assign t[167] = (x[56] & x[57]);
  assign t[168] = (x[20] & x[61]);
  assign t[169] = (x[34] & x[63]);
  assign t[16] = ~(t[114] & t[115]);
  assign t[170] = (x[34] & x[65]);
  assign t[171] = (x[39] & x[67]);
  assign t[172] = (x[39] & x[69]);
  assign t[173] = (x[71] & x[72]);
  assign t[174] = (x[25] & x[74]);
  assign t[175] = (x[48] & x[76]);
  assign t[176] = (x[48] & x[78]);
  assign t[177] = (x[51] & x[80]);
  assign t[178] = (x[51] & x[82]);
  assign t[179] = (x[84] & x[85]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[56] & x[87]);
  assign t[181] = (x[56] & x[89]);
  assign t[182] = (x[34] & x[91]);
  assign t[183] = (x[39] & x[93]);
  assign t[184] = (x[71] & x[95]);
  assign t[185] = (x[71] & x[97]);
  assign t[186] = (x[48] & x[99]);
  assign t[187] = (x[51] & x[101]);
  assign t[188] = (x[84] & x[103]);
  assign t[189] = (x[84] & x[105]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[56] & x[107]);
  assign t[191] = (x[71] & x[109]);
  assign t[192] = (x[84] & x[111]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[114]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[116]);
  assign t[31] = t[47] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = t[50] ^ t[42];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[54];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = ~(t[57] & t[117]);
  assign t[38] = t[58] ? x[29] : x[28];
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = t[63] ^ t[64];
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[40];
  assign t[44] = ~(t[118]);
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = ~(t[72] & t[120]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[17] ? x[38] : x[37];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[121]);
  assign t[53] = t[47] ? x[43] : x[42];
  assign t[54] = ~(t[76] & t[77]);
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = ~(t[24]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[82] & t[124]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = ~(t[85] & t[125]);
  assign t[63] = t[58] ? x[55] : x[54];
  assign t[64] = ~(t[86] & t[87]);
  assign t[65] = ~(t[88] & t[89]);
  assign t[66] = ~(t[90] & t[126]);
  assign t[67] = t[114] ? x[60] : x[59];
  assign t[68] = ~(t[119] & t[118]);
  assign t[69] = ~(t[127]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[91] & t[92]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[93] & t[94]);
  assign t[76] = ~(t[95] & t[96]);
  assign t[77] = ~(t[97] & t[132]);
  assign t[78] = ~(t[123] & t[122]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[98] & t[99]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[103]);
  assign t[87] = ~(t[104] & t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[140]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[105] & t[106]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[131] & t[130]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[144]);
  assign t[97] = ~(t[107] & t[108]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[111];
endmodule

module R1ind172(x, y);
 input [94:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[132] ^ x[29];
  assign t[101] = t[133] ^ x[31];
  assign t[102] = t[134] ^ x[35];
  assign t[103] = t[135] ^ x[38];
  assign t[104] = t[136] ^ x[40];
  assign t[105] = t[137] ^ x[45];
  assign t[106] = t[138] ^ x[47];
  assign t[107] = t[139] ^ x[51];
  assign t[108] = t[140] ^ x[54];
  assign t[109] = t[141] ^ x[56];
  assign t[10] = ~(x[3]);
  assign t[110] = t[142] ^ x[59];
  assign t[111] = t[143] ^ x[61];
  assign t[112] = t[144] ^ x[66];
  assign t[113] = t[145] ^ x[68];
  assign t[114] = t[146] ^ x[72];
  assign t[115] = t[147] ^ x[74];
  assign t[116] = t[148] ^ x[77];
  assign t[117] = t[149] ^ x[79];
  assign t[118] = t[150] ^ x[81];
  assign t[119] = t[151] ^ x[83];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[152] ^ x[85];
  assign t[121] = t[153] ^ x[88];
  assign t[122] = t[154] ^ x[90];
  assign t[123] = t[155] ^ x[92];
  assign t[124] = t[156] ^ x[94];
  assign t[125] = (x[0] & x[1]);
  assign t[126] = (x[8] & x[9]);
  assign t[127] = (x[11] & x[12]);
  assign t[128] = (x[14] & x[15]);
  assign t[129] = (x[17] & x[18]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & x[21]);
  assign t[131] = (x[20] & x[23]);
  assign t[132] = (x[27] & x[28]);
  assign t[133] = (x[27] & x[30]);
  assign t[134] = (x[20] & x[34]);
  assign t[135] = (x[36] & x[37]);
  assign t[136] = (x[36] & x[39]);
  assign t[137] = (x[43] & x[44]);
  assign t[138] = (x[43] & x[46]);
  assign t[139] = (x[27] & x[50]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[52] & x[53]);
  assign t[141] = (x[52] & x[55]);
  assign t[142] = (x[57] & x[58]);
  assign t[143] = (x[57] & x[60]);
  assign t[144] = (x[64] & x[65]);
  assign t[145] = (x[64] & x[67]);
  assign t[146] = (x[36] & x[71]);
  assign t[147] = (x[43] & x[73]);
  assign t[148] = (x[75] & x[76]);
  assign t[149] = (x[75] & x[78]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[52] & x[80]);
  assign t[151] = (x[57] & x[82]);
  assign t[152] = (x[64] & x[84]);
  assign t[153] = (x[86] & x[87]);
  assign t[154] = (x[86] & x[89]);
  assign t[155] = (x[75] & x[91]);
  assign t[156] = (x[86] & x[93]);
  assign t[15] = ~(t[94] & t[95]);
  assign t[16] = ~(t[96] & t[97]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[20];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[24] = ~(t[96]);
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = x[4] ? t[41] : t[40];
  assign t[28] = x[4] ? t[43] : t[42];
  assign t[29] = ~(t[98] & t[44]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = t[46] ? x[26] : x[25];
  assign t[32] = ~(t[47] & t[48]);
  assign t[33] = t[49] ^ t[40];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[53];
  assign t[36] = ~(t[100] & t[54]);
  assign t[37] = ~(t[101] & t[55]);
  assign t[38] = t[46] ? x[33] : x[32];
  assign t[39] = ~(t[56] & t[57]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = t[60] ^ t[42];
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[64];
  assign t[44] = ~(t[102]);
  assign t[45] = ~(t[102] & t[65]);
  assign t[46] = ~(t[24]);
  assign t[47] = ~(t[103] & t[66]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = t[68] ? x[42] : x[41];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = t[46] ? x[49] : x[48];
  assign t[53] = ~(t[71] & t[72]);
  assign t[54] = ~(t[107]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = ~(t[108] & t[74]);
  assign t[57] = ~(t[109] & t[75]);
  assign t[58] = ~(t[110] & t[76]);
  assign t[59] = ~(t[111] & t[77]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[68] ? x[63] : x[62];
  assign t[61] = ~(t[112] & t[78]);
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = t[17] ? x[70] : x[69];
  assign t[64] = ~(t[80] & t[81]);
  assign t[65] = ~(t[98]);
  assign t[66] = ~(t[114]);
  assign t[67] = ~(t[114] & t[82]);
  assign t[68] = ~(t[24]);
  assign t[69] = ~(t[115]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[117] & t[85]);
  assign t[73] = ~(t[100]);
  assign t[74] = ~(t[118]);
  assign t[75] = ~(t[118] & t[86]);
  assign t[76] = ~(t[119]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[123]);
  assign t[85] = ~(t[123] & t[91]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[124]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[124] & t[92]);
  assign t[91] = ~(t[116]);
  assign t[92] = ~(t[121]);
  assign t[93] = t[125] ^ x[2];
  assign t[94] = t[126] ^ x[10];
  assign t[95] = t[127] ^ x[13];
  assign t[96] = t[128] ^ x[16];
  assign t[97] = t[129] ^ x[19];
  assign t[98] = t[130] ^ x[22];
  assign t[99] = t[131] ^ x[24];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[93];
endmodule

module R1ind173(x, y);
 input [112:0] x;
 output y;

 wire [285:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[140] ? x[69] : x[68];
  assign t[101] = ~(t[141] & t[142]);
  assign t[102] = ~(t[226]);
  assign t[103] = ~(t[215] | t[216]);
  assign t[104] = ~(t[227]);
  assign t[105] = ~(t[228]);
  assign t[106] = ~(t[143] | t[144]);
  assign t[107] = ~(t[145] | t[146]);
  assign t[108] = ~(t[229]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[147] | t[148]);
  assign t[111] = ~(t[149] | t[150]);
  assign t[112] = ~(t[231] | t[151]);
  assign t[113] = t[29] ? x[84] : x[83];
  assign t[114] = ~(t[152] & t[153]);
  assign t[115] = ~(t[232]);
  assign t[116] = ~(t[233]);
  assign t[117] = ~(t[154] | t[155]);
  assign t[118] = t[29] ? x[90] : x[89];
  assign t[119] = ~(t[156] & t[157]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[158] & t[159]);
  assign t[121] = ~(t[160] & t[159]);
  assign t[122] = ~(x[4] & t[161]);
  assign t[123] = ~(t[162] & t[159]);
  assign t[124] = ~(t[160] & t[208]);
  assign t[125] = ~(t[80] | t[163]);
  assign t[126] = ~(t[80] | t[164]);
  assign t[127] = t[205] ? t[165] : t[123];
  assign t[128] = ~(t[78] | t[166]);
  assign t[129] = ~(t[167]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[80] | t[168]);
  assign t[131] = ~(t[234]);
  assign t[132] = ~(t[221] | t[222]);
  assign t[133] = ~(t[235]);
  assign t[134] = ~(t[236]);
  assign t[135] = ~(t[169] | t[170]);
  assign t[136] = ~(t[171] | t[126]);
  assign t[137] = ~(t[172] | t[173]);
  assign t[138] = ~(t[237]);
  assign t[139] = ~(t[224] | t[225]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[47]);
  assign t[141] = ~(t[174] | t[175]);
  assign t[142] = ~(t[176]);
  assign t[143] = ~(t[238]);
  assign t[144] = ~(t[227] | t[228]);
  assign t[145] = ~(t[30] & t[177]);
  assign t[146] = ~(t[178] & t[84]);
  assign t[147] = ~(t[239]);
  assign t[148] = ~(t[229] | t[230]);
  assign t[149] = ~(t[240]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[241]);
  assign t[151] = ~(t[179] | t[180]);
  assign t[152] = ~(t[125] | t[171]);
  assign t[153] = ~(t[181] | t[182]);
  assign t[154] = ~(t[242]);
  assign t[155] = ~(t[232] | t[233]);
  assign t[156] = ~(t[176] | t[50]);
  assign t[157] = ~(t[48] | t[183]);
  assign t[158] = x[4] & t[206];
  assign t[159] = ~(t[208]);
  assign t[15] = ~(t[205] & t[206]);
  assign t[160] = ~(x[4] | t[206]);
  assign t[161] = ~(t[206] | t[159]);
  assign t[162] = ~(x[4] | t[184]);
  assign t[163] = t[205] ? t[185] : t[121];
  assign t[164] = t[205] ? t[120] : t[124];
  assign t[165] = ~(x[4] & t[186]);
  assign t[166] = t[205] ? t[123] : t[165];
  assign t[167] = ~(t[174] | t[126]);
  assign t[168] = t[205] ? t[187] : t[165];
  assign t[169] = ~(t[243]);
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = ~(t[235] | t[236]);
  assign t[171] = ~(t[80] | t[188]);
  assign t[172] = t[208] & t[189];
  assign t[173] = ~(t[190]);
  assign t[174] = ~(t[80] | t[191]);
  assign t[175] = ~(t[192] & t[190]);
  assign t[176] = ~(t[80] | t[193]);
  assign t[177] = ~(t[78] & t[194]);
  assign t[178] = ~(t[172] & t[195]);
  assign t[179] = ~(t[244]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[240] | t[241]);
  assign t[181] = t[183] | t[130];
  assign t[182] = ~(t[196] & t[84]);
  assign t[183] = ~(t[190] & t[197]);
  assign t[184] = ~(t[206]);
  assign t[185] = ~(t[158] & t[208]);
  assign t[186] = ~(t[206] | t[208]);
  assign t[187] = ~(t[208] & t[162]);
  assign t[188] = t[205] ? t[165] : t[187];
  assign t[189] = ~(t[78] | t[205]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[198] | t[128]);
  assign t[191] = t[205] ? t[122] : t[123];
  assign t[192] = ~(t[125] | t[145]);
  assign t[193] = t[205] ? t[121] : t[185];
  assign t[194] = ~(t[165] & t[187]);
  assign t[195] = t[160] | t[158];
  assign t[196] = ~(t[199] | t[174]);
  assign t[197] = ~(t[161] & t[200]);
  assign t[198] = ~(t[78] | t[201]);
  assign t[199] = ~(t[202]);
  assign t[19] = t[29] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[80] & t[205];
  assign t[201] = t[205] ? t[120] : t[121];
  assign t[202] = ~(t[189] & t[203]);
  assign t[203] = ~(t[187] & t[122]);
  assign t[204] = t[245] ^ x[2];
  assign t[205] = t[246] ^ x[10];
  assign t[206] = t[247] ^ x[13];
  assign t[207] = t[248] ^ x[16];
  assign t[208] = t[249] ^ x[19];
  assign t[209] = t[250] ^ x[22];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[251] ^ x[25];
  assign t[211] = t[252] ^ x[27];
  assign t[212] = t[253] ^ x[29];
  assign t[213] = t[254] ^ x[34];
  assign t[214] = t[255] ^ x[37];
  assign t[215] = t[256] ^ x[39];
  assign t[216] = t[257] ^ x[41];
  assign t[217] = t[258] ^ x[44];
  assign t[218] = t[259] ^ x[49];
  assign t[219] = t[260] ^ x[52];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[261] ^ x[54];
  assign t[221] = t[262] ^ x[56];
  assign t[222] = t[263] ^ x[58];
  assign t[223] = t[264] ^ x[61];
  assign t[224] = t[265] ^ x[65];
  assign t[225] = t[266] ^ x[67];
  assign t[226] = t[267] ^ x[71];
  assign t[227] = t[268] ^ x[73];
  assign t[228] = t[269] ^ x[75];
  assign t[229] = t[270] ^ x[77];
  assign t[22] = ~(t[21] ^ t[34]);
  assign t[230] = t[271] ^ x[79];
  assign t[231] = t[272] ^ x[82];
  assign t[232] = t[273] ^ x[86];
  assign t[233] = t[274] ^ x[88];
  assign t[234] = t[275] ^ x[92];
  assign t[235] = t[276] ^ x[94];
  assign t[236] = t[277] ^ x[96];
  assign t[237] = t[278] ^ x[98];
  assign t[238] = t[279] ^ x[100];
  assign t[239] = t[280] ^ x[102];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[240] = t[281] ^ x[104];
  assign t[241] = t[282] ^ x[106];
  assign t[242] = t[283] ^ x[108];
  assign t[243] = t[284] ^ x[110];
  assign t[244] = t[285] ^ x[112];
  assign t[245] = (x[0] & x[1]);
  assign t[246] = (x[8] & x[9]);
  assign t[247] = (x[11] & x[12]);
  assign t[248] = (x[14] & x[15]);
  assign t[249] = (x[17] & x[18]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[20] & x[21]);
  assign t[251] = (x[23] & x[24]);
  assign t[252] = (x[20] & x[26]);
  assign t[253] = (x[20] & x[28]);
  assign t[254] = (x[32] & x[33]);
  assign t[255] = (x[35] & x[36]);
  assign t[256] = (x[23] & x[38]);
  assign t[257] = (x[23] & x[40]);
  assign t[258] = (x[42] & x[43]);
  assign t[259] = (x[47] & x[48]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[260] = (x[50] & x[51]);
  assign t[261] = (x[20] & x[53]);
  assign t[262] = (x[32] & x[55]);
  assign t[263] = (x[32] & x[57]);
  assign t[264] = (x[59] & x[60]);
  assign t[265] = (x[35] & x[64]);
  assign t[266] = (x[35] & x[66]);
  assign t[267] = (x[23] & x[70]);
  assign t[268] = (x[42] & x[72]);
  assign t[269] = (x[42] & x[74]);
  assign t[26] = ~(t[41] ^ t[42]);
  assign t[270] = (x[47] & x[76]);
  assign t[271] = (x[47] & x[78]);
  assign t[272] = (x[80] & x[81]);
  assign t[273] = (x[50] & x[85]);
  assign t[274] = (x[50] & x[87]);
  assign t[275] = (x[32] & x[91]);
  assign t[276] = (x[59] & x[93]);
  assign t[277] = (x[59] & x[95]);
  assign t[278] = (x[35] & x[97]);
  assign t[279] = (x[42] & x[99]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[280] = (x[47] & x[101]);
  assign t[281] = (x[80] & x[103]);
  assign t[282] = (x[80] & x[105]);
  assign t[283] = (x[50] & x[107]);
  assign t[284] = (x[59] & x[109]);
  assign t[285] = (x[80] & x[111]);
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[29] = ~(t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[209] | t[54]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[37] = ~(t[61] | t[62]);
  assign t[38] = ~(t[45] ^ t[63]);
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[210] | t[66]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[42] = ~(t[69] ^ t[70]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[45] = ~(t[75] | t[76]);
  assign t[46] = ~(t[43] ^ t[77]);
  assign t[47] = ~(t[207]);
  assign t[48] = ~(t[78] | t[79]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[80] | t[82]);
  assign t[51] = ~(t[83] & t[84]);
  assign t[52] = ~(t[211]);
  assign t[53] = ~(t[212]);
  assign t[54] = ~(t[85] | t[86]);
  assign t[55] = t[87] ? x[31] : x[30];
  assign t[56] = ~(t[88] & t[89]);
  assign t[57] = ~(t[90] | t[91]);
  assign t[58] = ~(t[213] | t[92]);
  assign t[59] = ~(t[93] | t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] ^ t[96]);
  assign t[61] = ~(t[97] | t[98]);
  assign t[62] = ~(t[214] | t[99]);
  assign t[63] = ~(t[100] ^ t[101]);
  assign t[64] = ~(t[215]);
  assign t[65] = ~(t[216]);
  assign t[66] = ~(t[102] | t[103]);
  assign t[67] = ~(t[104] | t[105]);
  assign t[68] = ~(t[217] | t[106]);
  assign t[69] = t[29] ? x[46] : x[45];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[107] & t[83]);
  assign t[71] = ~(t[108] | t[109]);
  assign t[72] = ~(t[218] | t[110]);
  assign t[73] = ~(t[111] | t[112]);
  assign t[74] = ~(t[113] ^ t[114]);
  assign t[75] = ~(t[115] | t[116]);
  assign t[76] = ~(t[219] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[207]);
  assign t[79] = t[205] ? t[121] : t[120];
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[78]);
  assign t[81] = t[205] ? t[123] : t[122];
  assign t[82] = t[205] ? t[124] : t[120];
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = t[78] | t[127];
  assign t[85] = ~(t[220]);
  assign t[86] = ~(t[211] | t[212]);
  assign t[87] = ~(t[47]);
  assign t[88] = ~(t[48] | t[128]);
  assign t[89] = ~(t[129] | t[130]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[221]);
  assign t[91] = ~(t[222]);
  assign t[92] = ~(t[131] | t[132]);
  assign t[93] = ~(t[133] | t[134]);
  assign t[94] = ~(t[223] | t[135]);
  assign t[95] = t[87] ? x[63] : x[62];
  assign t[96] = ~(t[136] & t[137]);
  assign t[97] = ~(t[224]);
  assign t[98] = ~(t[225]);
  assign t[99] = ~(t[138] | t[139]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[204];
endmodule

module R1ind174(x, y);
 input [121:0] x;
 output y;

 wire [198:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[107] | t[98]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[108] | t[103]);
  assign t[106] = ~(t[151]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = t[154] ^ x[2];
  assign t[10] = ~(x[3]);
  assign t[110] = t[155] ^ x[10];
  assign t[111] = t[156] ^ x[13];
  assign t[112] = t[157] ^ x[16];
  assign t[113] = t[158] ^ x[19];
  assign t[114] = t[159] ^ x[22];
  assign t[115] = t[160] ^ x[27];
  assign t[116] = t[161] ^ x[31];
  assign t[117] = t[162] ^ x[33];
  assign t[118] = t[163] ^ x[36];
  assign t[119] = t[164] ^ x[39];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[165] ^ x[44];
  assign t[121] = t[166] ^ x[48];
  assign t[122] = t[167] ^ x[50];
  assign t[123] = t[168] ^ x[53];
  assign t[124] = t[169] ^ x[56];
  assign t[125] = t[170] ^ x[61];
  assign t[126] = t[171] ^ x[65];
  assign t[127] = t[172] ^ x[67];
  assign t[128] = t[173] ^ x[69];
  assign t[129] = t[174] ^ x[71];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[73];
  assign t[131] = t[176] ^ x[75];
  assign t[132] = t[177] ^ x[77];
  assign t[133] = t[178] ^ x[80];
  assign t[134] = t[179] ^ x[82];
  assign t[135] = t[180] ^ x[84];
  assign t[136] = t[181] ^ x[86];
  assign t[137] = t[182] ^ x[88];
  assign t[138] = t[183] ^ x[90];
  assign t[139] = t[184] ^ x[93];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[95];
  assign t[141] = t[186] ^ x[97];
  assign t[142] = t[187] ^ x[99];
  assign t[143] = t[188] ^ x[101];
  assign t[144] = t[189] ^ x[103];
  assign t[145] = t[190] ^ x[105];
  assign t[146] = t[191] ^ x[107];
  assign t[147] = t[192] ^ x[109];
  assign t[148] = t[193] ^ x[111];
  assign t[149] = t[194] ^ x[113];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[115];
  assign t[151] = t[196] ^ x[117];
  assign t[152] = t[197] ^ x[119];
  assign t[153] = t[198] ^ x[121];
  assign t[154] = (x[0] & x[1]);
  assign t[155] = (x[8] & x[9]);
  assign t[156] = (x[11] & x[12]);
  assign t[157] = (x[14] & x[15]);
  assign t[158] = (x[17] & x[18]);
  assign t[159] = (x[20] & x[21]);
  assign t[15] = ~(t[110] & t[111]);
  assign t[160] = (x[25] & x[26]);
  assign t[161] = (x[20] & x[30]);
  assign t[162] = (x[20] & x[32]);
  assign t[163] = (x[34] & x[35]);
  assign t[164] = (x[37] & x[38]);
  assign t[165] = (x[42] & x[43]);
  assign t[166] = (x[25] & x[47]);
  assign t[167] = (x[25] & x[49]);
  assign t[168] = (x[51] & x[52]);
  assign t[169] = (x[54] & x[55]);
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = (x[59] & x[60]);
  assign t[171] = (x[20] & x[64]);
  assign t[172] = (x[34] & x[66]);
  assign t[173] = (x[34] & x[68]);
  assign t[174] = (x[37] & x[70]);
  assign t[175] = (x[37] & x[72]);
  assign t[176] = (x[42] & x[74]);
  assign t[177] = (x[42] & x[76]);
  assign t[178] = (x[78] & x[79]);
  assign t[179] = (x[25] & x[81]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[51] & x[83]);
  assign t[181] = (x[51] & x[85]);
  assign t[182] = (x[54] & x[87]);
  assign t[183] = (x[54] & x[89]);
  assign t[184] = (x[91] & x[92]);
  assign t[185] = (x[59] & x[94]);
  assign t[186] = (x[59] & x[96]);
  assign t[187] = (x[34] & x[98]);
  assign t[188] = (x[37] & x[100]);
  assign t[189] = (x[42] & x[102]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[78] & x[104]);
  assign t[191] = (x[78] & x[106]);
  assign t[192] = (x[51] & x[108]);
  assign t[193] = (x[54] & x[110]);
  assign t[194] = (x[91] & x[112]);
  assign t[195] = (x[91] & x[114]);
  assign t[196] = (x[59] & x[116]);
  assign t[197] = (x[78] & x[118]);
  assign t[198] = (x[91] & x[120]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[112]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[47] | t[114];
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[35];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[56];
  assign t[37] = ~(t[57] & t[58]);
  assign t[38] = t[59] | t[115];
  assign t[39] = t[60] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = t[69] ^ t[41];
  assign t[45] = ~(t[116]);
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[70] | t[45]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = t[73] | t[118];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = t[76] | t[119];
  assign t[52] = t[77] ? x[41] : x[40];
  assign t[53] = ~(t[78] & t[79]);
  assign t[54] = t[80] | t[120];
  assign t[55] = t[77] ? x[46] : x[45];
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = ~(t[121]);
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[83] | t[57]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[24]);
  assign t[61] = ~(t[84] & t[85]);
  assign t[62] = t[86] | t[123];
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = t[89] | t[124];
  assign t[65] = t[17] ? x[58] : x[57];
  assign t[66] = ~(t[90] & t[91]);
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = t[94] | t[125];
  assign t[69] = t[17] ? x[63] : x[62];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[95] | t[71]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[96] | t[74]);
  assign t[77] = ~(t[24]);
  assign t[78] = ~(t[131]);
  assign t[79] = ~(t[132]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[97] | t[78]);
  assign t[81] = ~(t[98] & t[99]);
  assign t[82] = t[100] | t[133];
  assign t[83] = ~(t[134]);
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[101] | t[84]);
  assign t[87] = ~(t[137]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[102] | t[87]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[103] & t[104]);
  assign t[91] = t[105] | t[139];
  assign t[92] = ~(t[140]);
  assign t[93] = ~(t[141]);
  assign t[94] = ~(t[106] | t[92]);
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[109];
endmodule

module R1ind175(x, y);
 input [121:0] x;
 output y;

 wire [207:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[155]);
  assign t[104] = ~(t[114] & t[115]);
  assign t[105] = ~(t[145] & t[144]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[147] & t[146]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[159]);
  assign t[111] = ~(t[116] & t[117]);
  assign t[112] = ~(t[150] & t[149]);
  assign t[113] = ~(t[160]);
  assign t[114] = ~(t[155] & t[154]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[159] & t[158]);
  assign t[117] = ~(t[162]);
  assign t[118] = t[163] ^ x[2];
  assign t[119] = t[164] ^ x[10];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[165] ^ x[13];
  assign t[121] = t[166] ^ x[16];
  assign t[122] = t[167] ^ x[19];
  assign t[123] = t[168] ^ x[22];
  assign t[124] = t[169] ^ x[27];
  assign t[125] = t[170] ^ x[31];
  assign t[126] = t[171] ^ x[33];
  assign t[127] = t[172] ^ x[36];
  assign t[128] = t[173] ^ x[39];
  assign t[129] = t[174] ^ x[44];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[175] ^ x[48];
  assign t[131] = t[176] ^ x[50];
  assign t[132] = t[177] ^ x[53];
  assign t[133] = t[178] ^ x[56];
  assign t[134] = t[179] ^ x[61];
  assign t[135] = t[180] ^ x[65];
  assign t[136] = t[181] ^ x[67];
  assign t[137] = t[182] ^ x[69];
  assign t[138] = t[183] ^ x[71];
  assign t[139] = t[184] ^ x[73];
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = t[185] ^ x[75];
  assign t[141] = t[186] ^ x[77];
  assign t[142] = t[187] ^ x[80];
  assign t[143] = t[188] ^ x[82];
  assign t[144] = t[189] ^ x[84];
  assign t[145] = t[190] ^ x[86];
  assign t[146] = t[191] ^ x[88];
  assign t[147] = t[192] ^ x[90];
  assign t[148] = t[193] ^ x[93];
  assign t[149] = t[194] ^ x[95];
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = t[195] ^ x[97];
  assign t[151] = t[196] ^ x[99];
  assign t[152] = t[197] ^ x[101];
  assign t[153] = t[198] ^ x[103];
  assign t[154] = t[199] ^ x[105];
  assign t[155] = t[200] ^ x[107];
  assign t[156] = t[201] ^ x[109];
  assign t[157] = t[202] ^ x[111];
  assign t[158] = t[203] ^ x[113];
  assign t[159] = t[204] ^ x[115];
  assign t[15] = ~(t[119] & t[120]);
  assign t[160] = t[205] ^ x[117];
  assign t[161] = t[206] ^ x[119];
  assign t[162] = t[207] ^ x[121];
  assign t[163] = (x[0] & x[1]);
  assign t[164] = (x[8] & x[9]);
  assign t[165] = (x[11] & x[12]);
  assign t[166] = (x[14] & x[15]);
  assign t[167] = (x[17] & x[18]);
  assign t[168] = (x[20] & x[21]);
  assign t[169] = (x[25] & x[26]);
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = (x[20] & x[30]);
  assign t[171] = (x[20] & x[32]);
  assign t[172] = (x[34] & x[35]);
  assign t[173] = (x[37] & x[38]);
  assign t[174] = (x[42] & x[43]);
  assign t[175] = (x[25] & x[47]);
  assign t[176] = (x[25] & x[49]);
  assign t[177] = (x[51] & x[52]);
  assign t[178] = (x[54] & x[55]);
  assign t[179] = (x[59] & x[60]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[20] & x[64]);
  assign t[181] = (x[34] & x[66]);
  assign t[182] = (x[34] & x[68]);
  assign t[183] = (x[37] & x[70]);
  assign t[184] = (x[37] & x[72]);
  assign t[185] = (x[42] & x[74]);
  assign t[186] = (x[42] & x[76]);
  assign t[187] = (x[78] & x[79]);
  assign t[188] = (x[25] & x[81]);
  assign t[189] = (x[51] & x[83]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[190] = (x[51] & x[85]);
  assign t[191] = (x[54] & x[87]);
  assign t[192] = (x[54] & x[89]);
  assign t[193] = (x[91] & x[92]);
  assign t[194] = (x[59] & x[94]);
  assign t[195] = (x[59] & x[96]);
  assign t[196] = (x[34] & x[98]);
  assign t[197] = (x[37] & x[100]);
  assign t[198] = (x[42] & x[102]);
  assign t[199] = (x[78] & x[104]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = (x[78] & x[106]);
  assign t[201] = (x[51] & x[108]);
  assign t[202] = (x[54] & x[110]);
  assign t[203] = (x[91] & x[112]);
  assign t[204] = (x[91] & x[114]);
  assign t[205] = (x[59] & x[116]);
  assign t[206] = (x[78] & x[118]);
  assign t[207] = (x[91] & x[120]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[121]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[47] & t[123]);
  assign t[31] = t[17] ? x[24] : x[23];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[35];
  assign t[35] = ~(t[53] & t[54]);
  assign t[36] = t[55] ^ t[56];
  assign t[37] = ~(t[57] & t[58]);
  assign t[38] = ~(t[59] & t[124]);
  assign t[39] = t[60] ? x[29] : x[28];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = t[65] ^ t[66];
  assign t[43] = ~(t[67] & t[68]);
  assign t[44] = t[69] ^ t[41];
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = ~(t[74] & t[127]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[75] & t[76]);
  assign t[51] = ~(t[77] & t[128]);
  assign t[52] = t[60] ? x[41] : x[40];
  assign t[53] = ~(t[78] & t[79]);
  assign t[54] = ~(t[80] & t[129]);
  assign t[55] = t[60] ? x[46] : x[45];
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = ~(t[130]);
  assign t[58] = ~(t[131]);
  assign t[59] = ~(t[83] & t[84]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[24]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[87] & t[132]);
  assign t[63] = ~(t[88] & t[89]);
  assign t[64] = ~(t[90] & t[133]);
  assign t[65] = t[17] ? x[58] : x[57];
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = ~(t[93] & t[94]);
  assign t[68] = ~(t[95] & t[134]);
  assign t[69] = t[121] ? x[63] : x[62];
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[126] & t[125]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[96] & t[97]);
  assign t[75] = ~(t[138]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[98] & t[99]);
  assign t[78] = ~(t[140]);
  assign t[79] = ~(t[141]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[100] & t[101]);
  assign t[81] = ~(t[102] & t[103]);
  assign t[82] = ~(t[104] & t[142]);
  assign t[83] = ~(t[131] & t[130]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[105] & t[106]);
  assign t[88] = ~(t[146]);
  assign t[89] = ~(t[147]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[107] & t[108]);
  assign t[91] = ~(t[109] & t[110]);
  assign t[92] = ~(t[111] & t[148]);
  assign t[93] = ~(t[149]);
  assign t[94] = ~(t[150]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[118];
endmodule

module R1ind176(x, y);
 input [101:0] x;
 output y;

 wire [168:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[135] ^ x[10];
  assign t[101] = t[136] ^ x[13];
  assign t[102] = t[137] ^ x[16];
  assign t[103] = t[138] ^ x[19];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[24];
  assign t[106] = t[141] ^ x[29];
  assign t[107] = t[142] ^ x[31];
  assign t[108] = t[143] ^ x[35];
  assign t[109] = t[144] ^ x[38];
  assign t[10] = ~(x[3]);
  assign t[110] = t[145] ^ x[40];
  assign t[111] = t[146] ^ x[43];
  assign t[112] = t[147] ^ x[45];
  assign t[113] = t[148] ^ x[50];
  assign t[114] = t[149] ^ x[52];
  assign t[115] = t[150] ^ x[56];
  assign t[116] = t[151] ^ x[59];
  assign t[117] = t[152] ^ x[61];
  assign t[118] = t[153] ^ x[64];
  assign t[119] = t[154] ^ x[66];
  assign t[11] = t[17] ? x[6] : x[7];
  assign t[120] = t[155] ^ x[71];
  assign t[121] = t[156] ^ x[73];
  assign t[122] = t[157] ^ x[77];
  assign t[123] = t[158] ^ x[79];
  assign t[124] = t[159] ^ x[82];
  assign t[125] = t[160] ^ x[84];
  assign t[126] = t[161] ^ x[86];
  assign t[127] = t[162] ^ x[88];
  assign t[128] = t[163] ^ x[90];
  assign t[129] = t[164] ^ x[92];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[165] ^ x[95];
  assign t[131] = t[166] ^ x[97];
  assign t[132] = t[167] ^ x[99];
  assign t[133] = t[168] ^ x[101];
  assign t[134] = (x[0] & x[1]);
  assign t[135] = (x[8] & x[9]);
  assign t[136] = (x[11] & x[12]);
  assign t[137] = (x[14] & x[15]);
  assign t[138] = (x[17] & x[18]);
  assign t[139] = (x[20] & x[21]);
  assign t[13] = x[4] ? t[21] : t[20];
  assign t[140] = (x[20] & x[23]);
  assign t[141] = (x[27] & x[28]);
  assign t[142] = (x[27] & x[30]);
  assign t[143] = (x[20] & x[34]);
  assign t[144] = (x[36] & x[37]);
  assign t[145] = (x[36] & x[39]);
  assign t[146] = (x[41] & x[42]);
  assign t[147] = (x[41] & x[44]);
  assign t[148] = (x[48] & x[49]);
  assign t[149] = (x[48] & x[51]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[150] = (x[27] & x[55]);
  assign t[151] = (x[57] & x[58]);
  assign t[152] = (x[57] & x[60]);
  assign t[153] = (x[62] & x[63]);
  assign t[154] = (x[62] & x[65]);
  assign t[155] = (x[69] & x[70]);
  assign t[156] = (x[69] & x[72]);
  assign t[157] = (x[36] & x[76]);
  assign t[158] = (x[41] & x[78]);
  assign t[159] = (x[80] & x[81]);
  assign t[15] = ~(t[100] & t[101]);
  assign t[160] = (x[80] & x[83]);
  assign t[161] = (x[48] & x[85]);
  assign t[162] = (x[57] & x[87]);
  assign t[163] = (x[62] & x[89]);
  assign t[164] = (x[69] & x[91]);
  assign t[165] = (x[93] & x[94]);
  assign t[166] = (x[93] & x[96]);
  assign t[167] = (x[80] & x[98]);
  assign t[168] = (x[93] & x[100]);
  assign t[16] = ~(t[102] & t[103]);
  assign t[17] = ~(t[24]);
  assign t[18] = x[4] ? t[26] : t[25];
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = t[31] ^ t[32];
  assign t[22] = x[4] ? t[34] : t[33];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[24] = ~(t[102]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[39] ^ t[40];
  assign t[27] = x[4] ? t[42] : t[41];
  assign t[28] = x[4] ? t[44] : t[43];
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = t[47] ? x[26] : x[25];
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = t[56] ^ t[33];
  assign t[37] = ~(t[106] & t[57]);
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = t[47] ? x[33] : x[32];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[43];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[108]);
  assign t[46] = ~(t[108] & t[68]);
  assign t[47] = ~(t[24]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = t[73] ? x[47] : x[46];
  assign t[53] = ~(t[74] & t[75]);
  assign t[54] = ~(t[113] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = t[73] ? x[54] : x[53];
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = t[73] ? x[68] : x[67];
  assign t[64] = ~(t[120] & t[83]);
  assign t[65] = ~(t[121] & t[84]);
  assign t[66] = t[47] ? x[75] : x[74];
  assign t[67] = ~(t[85] & t[86]);
  assign t[68] = ~(t[104]);
  assign t[69] = ~(t[122]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[122] & t[87]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[24]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126]);
  assign t[77] = ~(t[126] & t[91]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[127]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[127] & t[92]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[132]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[132] & t[97]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[118]);
  assign t[94] = ~(t[120]);
  assign t[95] = ~(t[133]);
  assign t[96] = ~(t[133] & t[98]);
  assign t[97] = ~(t[124]);
  assign t[98] = ~(t[130]);
  assign t[99] = t[134] ^ x[2];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind177(x, y);
 input [121:0] x;
 output y;

 wire [293:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[226]);
  assign t[101] = ~(t[227]);
  assign t[102] = ~(t[145] | t[146]);
  assign t[103] = ~(t[147] | t[148]);
  assign t[104] = ~(t[228] | t[149]);
  assign t[105] = t[142] ? x[76] : x[75];
  assign t[106] = ~(t[150] & t[151]);
  assign t[107] = ~(t[229]);
  assign t[108] = ~(t[216] | t[217]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[152] | t[153]);
  assign t[112] = ~(t[154] | t[155]);
  assign t[113] = ~(t[232]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[156] | t[157]);
  assign t[116] = ~(t[158] | t[159]);
  assign t[117] = ~(t[234] | t[160]);
  assign t[118] = t[29] ? x[91] : x[90];
  assign t[119] = ~(t[161] & t[162]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[235]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[163] | t[164]);
  assign t[123] = t[29] ? x[97] : x[96];
  assign t[124] = ~(t[165] & t[166]);
  assign t[125] = ~(t[127] | t[167]);
  assign t[126] = ~(t[85] | t[168]);
  assign t[127] = ~(t[207]);
  assign t[128] = ~(t[169] & t[170]);
  assign t[129] = t[208] & t[171];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = t[172] | t[173];
  assign t[131] = t[205] ? t[169] : t[174];
  assign t[132] = ~(t[172] & t[175]);
  assign t[133] = ~(t[173] & t[208]);
  assign t[134] = ~(t[172] & t[208]);
  assign t[135] = ~(t[173] & t[175]);
  assign t[136] = ~(t[237]);
  assign t[137] = ~(t[222] | t[223]);
  assign t[138] = ~(t[206] | t[175]);
  assign t[139] = t[85] & t[205];
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[238]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[48]);
  assign t[143] = ~(t[176] & t[94]);
  assign t[144] = ~(t[85] | t[177]);
  assign t[145] = ~(t[239]);
  assign t[146] = ~(t[226] | t[227]);
  assign t[147] = ~(t[240]);
  assign t[148] = ~(t[241]);
  assign t[149] = ~(t[178] | t[179]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[51]);
  assign t[151] = ~(t[180] | t[144]);
  assign t[152] = ~(t[242]);
  assign t[153] = ~(t[230] | t[231]);
  assign t[154] = ~(t[85] | t[181]);
  assign t[155] = ~(t[31] & t[84]);
  assign t[156] = ~(t[243]);
  assign t[157] = ~(t[232] | t[233]);
  assign t[158] = ~(t[244]);
  assign t[159] = ~(t[245]);
  assign t[15] = ~(t[205] & t[206]);
  assign t[160] = ~(t[182] | t[183]);
  assign t[161] = ~(t[51] | t[184]);
  assign t[162] = ~(t[99] | t[185]);
  assign t[163] = ~(t[246]);
  assign t[164] = ~(t[235] | t[236]);
  assign t[165] = ~(t[186] | t[154]);
  assign t[166] = ~(t[125] | t[143]);
  assign t[167] = t[205] ? t[132] : t[135];
  assign t[168] = t[205] ? t[174] : t[187];
  assign t[169] = ~(x[4] & t[188]);
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = ~(t[208] & t[189]);
  assign t[171] = ~(t[127] | t[205]);
  assign t[172] = ~(x[4] | t[206]);
  assign t[173] = x[4] & t[206];
  assign t[174] = ~(t[189] & t[175]);
  assign t[175] = ~(t[208]);
  assign t[176] = ~(t[190] | t[191]);
  assign t[177] = t[205] ? t[170] : t[169];
  assign t[178] = ~(t[247]);
  assign t[179] = ~(t[240] | t[241]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[192]);
  assign t[181] = t[205] ? t[134] : t[135];
  assign t[182] = ~(t[248]);
  assign t[183] = ~(t[244] | t[245]);
  assign t[184] = ~(t[85] | t[193]);
  assign t[185] = ~(t[194] & t[84]);
  assign t[186] = ~(t[85] | t[195]);
  assign t[187] = ~(x[4] & t[138]);
  assign t[188] = ~(t[206] | t[208]);
  assign t[189] = ~(x[4] | t[196]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[127] | t[197]);
  assign t[191] = ~(t[127] | t[198]);
  assign t[192] = ~(t[199] | t[52]);
  assign t[193] = t[205] ? t[169] : t[170];
  assign t[194] = ~(t[200] | t[199]);
  assign t[195] = t[205] ? t[132] : t[133];
  assign t[196] = ~(t[206]);
  assign t[197] = t[205] ? t[135] : t[132];
  assign t[198] = t[205] ? t[174] : t[169];
  assign t[199] = ~(t[85] | t[201]);
  assign t[19] = t[29] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = ~(t[202]);
  assign t[201] = t[205] ? t[187] : t[174];
  assign t[202] = ~(t[171] & t[203]);
  assign t[203] = ~(t[170] & t[187]);
  assign t[204] = t[249] ^ x[2];
  assign t[205] = t[250] ^ x[10];
  assign t[206] = t[251] ^ x[13];
  assign t[207] = t[252] ^ x[16];
  assign t[208] = t[253] ^ x[19];
  assign t[209] = t[254] ^ x[22];
  assign t[20] = ~(t[30] & t[31]);
  assign t[210] = t[255] ^ x[25];
  assign t[211] = t[256] ^ x[27];
  assign t[212] = t[257] ^ x[29];
  assign t[213] = t[258] ^ x[32];
  assign t[214] = t[259] ^ x[37];
  assign t[215] = t[260] ^ x[40];
  assign t[216] = t[261] ^ x[42];
  assign t[217] = t[262] ^ x[44];
  assign t[218] = t[263] ^ x[47];
  assign t[219] = t[264] ^ x[52];
  assign t[21] = ~(t[32] | t[33]);
  assign t[220] = t[265] ^ x[55];
  assign t[221] = t[266] ^ x[57];
  assign t[222] = t[267] ^ x[59];
  assign t[223] = t[268] ^ x[61];
  assign t[224] = t[269] ^ x[63];
  assign t[225] = t[270] ^ x[65];
  assign t[226] = t[271] ^ x[69];
  assign t[227] = t[272] ^ x[71];
  assign t[228] = t[273] ^ x[74];
  assign t[229] = t[274] ^ x[78];
  assign t[22] = ~(t[34] ^ t[35]);
  assign t[230] = t[275] ^ x[80];
  assign t[231] = t[276] ^ x[82];
  assign t[232] = t[277] ^ x[84];
  assign t[233] = t[278] ^ x[86];
  assign t[234] = t[279] ^ x[89];
  assign t[235] = t[280] ^ x[93];
  assign t[236] = t[281] ^ x[95];
  assign t[237] = t[282] ^ x[99];
  assign t[238] = t[283] ^ x[101];
  assign t[239] = t[284] ^ x[103];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[240] = t[285] ^ x[105];
  assign t[241] = t[286] ^ x[107];
  assign t[242] = t[287] ^ x[109];
  assign t[243] = t[288] ^ x[111];
  assign t[244] = t[289] ^ x[113];
  assign t[245] = t[290] ^ x[115];
  assign t[246] = t[291] ^ x[117];
  assign t[247] = t[292] ^ x[119];
  assign t[248] = t[293] ^ x[121];
  assign t[249] = (x[0] & x[1]);
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[250] = (x[8] & x[9]);
  assign t[251] = (x[11] & x[12]);
  assign t[252] = (x[14] & x[15]);
  assign t[253] = (x[17] & x[18]);
  assign t[254] = (x[20] & x[21]);
  assign t[255] = (x[23] & x[24]);
  assign t[256] = (x[20] & x[26]);
  assign t[257] = (x[20] & x[28]);
  assign t[258] = (x[30] & x[31]);
  assign t[259] = (x[35] & x[36]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[260] = (x[38] & x[39]);
  assign t[261] = (x[23] & x[41]);
  assign t[262] = (x[23] & x[43]);
  assign t[263] = (x[45] & x[46]);
  assign t[264] = (x[50] & x[51]);
  assign t[265] = (x[53] & x[54]);
  assign t[266] = (x[20] & x[56]);
  assign t[267] = (x[30] & x[58]);
  assign t[268] = (x[30] & x[60]);
  assign t[269] = (x[35] & x[62]);
  assign t[26] = ~(t[42] ^ t[43]);
  assign t[270] = (x[35] & x[64]);
  assign t[271] = (x[38] & x[68]);
  assign t[272] = (x[38] & x[70]);
  assign t[273] = (x[72] & x[73]);
  assign t[274] = (x[23] & x[77]);
  assign t[275] = (x[45] & x[79]);
  assign t[276] = (x[45] & x[81]);
  assign t[277] = (x[50] & x[83]);
  assign t[278] = (x[50] & x[85]);
  assign t[279] = (x[87] & x[88]);
  assign t[27] = x[4] ? t[45] : t[44];
  assign t[280] = (x[53] & x[92]);
  assign t[281] = (x[53] & x[94]);
  assign t[282] = (x[30] & x[98]);
  assign t[283] = (x[35] & x[100]);
  assign t[284] = (x[38] & x[102]);
  assign t[285] = (x[72] & x[104]);
  assign t[286] = (x[72] & x[106]);
  assign t[287] = (x[45] & x[108]);
  assign t[288] = (x[50] & x[110]);
  assign t[289] = (x[87] & x[112]);
  assign t[28] = x[4] ? t[47] : t[46];
  assign t[290] = (x[87] & x[114]);
  assign t[291] = (x[53] & x[116]);
  assign t[292] = (x[72] & x[118]);
  assign t[293] = (x[87] & x[120]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51] | t[52]);
  assign t[32] = ~(t[53] | t[54]);
  assign t[33] = ~(t[209] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[58] ^ t[59]);
  assign t[36] = ~(t[60] | t[61]);
  assign t[37] = ~(t[38] ^ t[62]);
  assign t[38] = ~(t[63] | t[64]);
  assign t[39] = ~(t[65] ^ t[66]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[67] | t[68]);
  assign t[41] = ~(t[210] | t[69]);
  assign t[42] = ~(t[70] | t[71]);
  assign t[43] = ~(t[72] ^ t[73]);
  assign t[44] = ~(t[74] | t[75]);
  assign t[45] = ~(t[76] ^ t[77]);
  assign t[46] = ~(t[78] | t[79]);
  assign t[47] = ~(t[44] ^ t[80]);
  assign t[48] = ~(t[207]);
  assign t[49] = ~(t[81] & t[82]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[83] & t[84]);
  assign t[51] = ~(t[85] | t[86]);
  assign t[52] = ~(t[85] | t[87]);
  assign t[53] = ~(t[211]);
  assign t[54] = ~(t[212]);
  assign t[55] = ~(t[88] | t[89]);
  assign t[56] = ~(t[90] | t[91]);
  assign t[57] = ~(t[213] | t[92]);
  assign t[58] = t[29] ? x[34] : x[33];
  assign t[59] = ~(t[93] & t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[214] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[100] | t[101]);
  assign t[64] = ~(t[215] | t[102]);
  assign t[65] = ~(t[103] | t[104]);
  assign t[66] = ~(t[105] ^ t[106]);
  assign t[67] = ~(t[216]);
  assign t[68] = ~(t[217]);
  assign t[69] = ~(t[107] | t[108]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[109] | t[110]);
  assign t[71] = ~(t[218] | t[111]);
  assign t[72] = t[29] ? x[49] : x[48];
  assign t[73] = ~(t[81] & t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[219] | t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[120] | t[121]);
  assign t[79] = ~(t[220] | t[122]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[123] ^ t[124]);
  assign t[81] = ~(t[125] | t[126]);
  assign t[82] = ~(t[127] & t[128]);
  assign t[83] = ~(t[129] & t[130]);
  assign t[84] = t[127] | t[131];
  assign t[85] = ~(t[127]);
  assign t[86] = t[205] ? t[133] : t[132];
  assign t[87] = t[205] ? t[135] : t[134];
  assign t[88] = ~(t[221]);
  assign t[89] = ~(t[211] | t[212]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[222]);
  assign t[91] = ~(t[223]);
  assign t[92] = ~(t[136] | t[137]);
  assign t[93] = ~(t[51] | t[49]);
  assign t[94] = ~(t[138] & t[139]);
  assign t[95] = ~(t[224]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[140] | t[141]);
  assign t[98] = t[142] ? x[67] : x[66];
  assign t[99] = t[143] | t[144];
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[204];
endmodule

module R1ind178(x, y);
 input [112:0] x;
 output y;

 wire [180:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[141] ^ x[8];
  assign t[101] = t[142] ^ x[11];
  assign t[102] = t[143] ^ x[14];
  assign t[103] = t[144] ^ x[17];
  assign t[104] = t[145] ^ x[22];
  assign t[105] = t[146] ^ x[27];
  assign t[106] = t[147] ^ x[31];
  assign t[107] = t[148] ^ x[33];
  assign t[108] = t[149] ^ x[36];
  assign t[109] = t[150] ^ x[39];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[151] ^ x[44];
  assign t[111] = t[152] ^ x[48];
  assign t[112] = t[153] ^ x[50];
  assign t[113] = t[154] ^ x[53];
  assign t[114] = t[155] ^ x[58];
  assign t[115] = t[156] ^ x[62];
  assign t[116] = t[157] ^ x[64];
  assign t[117] = t[158] ^ x[66];
  assign t[118] = t[159] ^ x[68];
  assign t[119] = t[160] ^ x[70];
  assign t[11] = t[102] ? x[18] : x[19];
  assign t[120] = t[161] ^ x[72];
  assign t[121] = t[162] ^ x[74];
  assign t[122] = t[163] ^ x[76];
  assign t[123] = t[164] ^ x[78];
  assign t[124] = t[165] ^ x[80];
  assign t[125] = t[166] ^ x[83];
  assign t[126] = t[167] ^ x[85];
  assign t[127] = t[168] ^ x[87];
  assign t[128] = t[169] ^ x[90];
  assign t[129] = t[170] ^ x[92];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = t[171] ^ x[94];
  assign t[131] = t[172] ^ x[96];
  assign t[132] = t[173] ^ x[98];
  assign t[133] = t[174] ^ x[100];
  assign t[134] = t[175] ^ x[102];
  assign t[135] = t[176] ^ x[104];
  assign t[136] = t[177] ^ x[106];
  assign t[137] = t[178] ^ x[108];
  assign t[138] = t[179] ^ x[110];
  assign t[139] = t[180] ^ x[112];
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (x[0] & x[1]);
  assign t[141] = (x[6] & x[7]);
  assign t[142] = (x[9] & x[10]);
  assign t[143] = (x[12] & x[13]);
  assign t[144] = (x[15] & x[16]);
  assign t[145] = (x[20] & x[21]);
  assign t[146] = (x[25] & x[26]);
  assign t[147] = (x[20] & x[30]);
  assign t[148] = (x[20] & x[32]);
  assign t[149] = (x[34] & x[35]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[37] & x[38]);
  assign t[151] = (x[42] & x[43]);
  assign t[152] = (x[25] & x[47]);
  assign t[153] = (x[25] & x[49]);
  assign t[154] = (x[51] & x[52]);
  assign t[155] = (x[56] & x[57]);
  assign t[156] = (x[20] & x[61]);
  assign t[157] = (x[34] & x[63]);
  assign t[158] = (x[34] & x[65]);
  assign t[159] = (x[37] & x[67]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[160] = (x[37] & x[69]);
  assign t[161] = (x[42] & x[71]);
  assign t[162] = (x[42] & x[73]);
  assign t[163] = (x[25] & x[75]);
  assign t[164] = (x[51] & x[77]);
  assign t[165] = (x[51] & x[79]);
  assign t[166] = (x[81] & x[82]);
  assign t[167] = (x[56] & x[84]);
  assign t[168] = (x[56] & x[86]);
  assign t[169] = (x[88] & x[89]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (x[34] & x[91]);
  assign t[171] = (x[37] & x[93]);
  assign t[172] = (x[42] & x[95]);
  assign t[173] = (x[51] & x[97]);
  assign t[174] = (x[81] & x[99]);
  assign t[175] = (x[81] & x[101]);
  assign t[176] = (x[56] & x[103]);
  assign t[177] = (x[88] & x[105]);
  assign t[178] = (x[88] & x[107]);
  assign t[179] = (x[81] & x[109]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[180] = (x[88] & x[111]);
  assign t[18] = t[27] ^ t[28];
  assign t[19] = x[4] ? t[30] : t[29];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = t[35] ^ t[21];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[40] & t[41]);
  assign t[26] = t[42] | t[104];
  assign t[27] = t[43] ? x[24] : x[23];
  assign t[28] = ~(t[44] & t[45]);
  assign t[29] = ~(t[46] & t[47]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[48] ^ t[36];
  assign t[31] = ~(t[49] & t[50]);
  assign t[32] = t[51] ^ t[29];
  assign t[33] = ~(t[52] & t[53]);
  assign t[34] = t[54] | t[105];
  assign t[35] = t[102] ? x[29] : x[28];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[58];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[106]);
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[63] | t[40]);
  assign t[43] = ~(t[64]);
  assign t[44] = ~(t[65] & t[66]);
  assign t[45] = t[67] | t[108];
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = t[70] | t[109];
  assign t[48] = t[43] ? x[41] : x[40];
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[73] | t[110];
  assign t[51] = t[43] ? x[46] : x[45];
  assign t[52] = ~(t[111]);
  assign t[53] = ~(t[112]);
  assign t[54] = ~(t[74] | t[52]);
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = t[77] | t[113];
  assign t[57] = t[102] ? x[55] : x[54];
  assign t[58] = ~(t[78] & t[79]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = t[82] | t[114];
  assign t[61] = t[83] ? x[60] : x[59];
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = ~(t[115]);
  assign t[64] = ~(t[102]);
  assign t[65] = ~(t[116]);
  assign t[66] = ~(t[117]);
  assign t[67] = ~(t[86] | t[65]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[119]);
  assign t[6] = ~(t[100] & t[101]);
  assign t[70] = ~(t[87] | t[68]);
  assign t[71] = ~(t[120]);
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[88] | t[71]);
  assign t[74] = ~(t[122]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[89] | t[75]);
  assign t[78] = ~(t[90] & t[91]);
  assign t[79] = t[92] | t[125];
  assign t[7] = ~(t[102] & t[103]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[93] | t[80]);
  assign t[83] = ~(t[64]);
  assign t[84] = ~(t[94] & t[95]);
  assign t[85] = t[96] | t[128];
  assign t[86] = ~(t[129]);
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[97] | t[90]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[98] | t[94]);
  assign t[97] = ~(t[138]);
  assign t[98] = ~(t[139]);
  assign t[99] = t[140] ^ x[2];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind179(x, y);
 input [112:0] x;
 output y;

 wire [188:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[144]);
  assign t[101] = ~(t[145]);
  assign t[102] = ~(t[105] & t[106]);
  assign t[103] = ~(t[142] & t[141]);
  assign t[104] = ~(t[146]);
  assign t[105] = ~(t[145] & t[144]);
  assign t[106] = ~(t[147]);
  assign t[107] = t[148] ^ x[2];
  assign t[108] = t[149] ^ x[8];
  assign t[109] = t[150] ^ x[11];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[151] ^ x[14];
  assign t[111] = t[152] ^ x[17];
  assign t[112] = t[153] ^ x[22];
  assign t[113] = t[154] ^ x[27];
  assign t[114] = t[155] ^ x[31];
  assign t[115] = t[156] ^ x[33];
  assign t[116] = t[157] ^ x[36];
  assign t[117] = t[158] ^ x[39];
  assign t[118] = t[159] ^ x[44];
  assign t[119] = t[160] ^ x[48];
  assign t[11] = t[110] ? x[18] : x[19];
  assign t[120] = t[161] ^ x[50];
  assign t[121] = t[162] ^ x[53];
  assign t[122] = t[163] ^ x[58];
  assign t[123] = t[164] ^ x[62];
  assign t[124] = t[165] ^ x[64];
  assign t[125] = t[166] ^ x[66];
  assign t[126] = t[167] ^ x[68];
  assign t[127] = t[168] ^ x[70];
  assign t[128] = t[169] ^ x[72];
  assign t[129] = t[170] ^ x[74];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = t[171] ^ x[76];
  assign t[131] = t[172] ^ x[78];
  assign t[132] = t[173] ^ x[80];
  assign t[133] = t[174] ^ x[83];
  assign t[134] = t[175] ^ x[85];
  assign t[135] = t[176] ^ x[87];
  assign t[136] = t[177] ^ x[90];
  assign t[137] = t[178] ^ x[92];
  assign t[138] = t[179] ^ x[94];
  assign t[139] = t[180] ^ x[96];
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = t[181] ^ x[98];
  assign t[141] = t[182] ^ x[100];
  assign t[142] = t[183] ^ x[102];
  assign t[143] = t[184] ^ x[104];
  assign t[144] = t[185] ^ x[106];
  assign t[145] = t[186] ^ x[108];
  assign t[146] = t[187] ^ x[110];
  assign t[147] = t[188] ^ x[112];
  assign t[148] = (x[0] & x[1]);
  assign t[149] = (x[6] & x[7]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[9] & x[10]);
  assign t[151] = (x[12] & x[13]);
  assign t[152] = (x[15] & x[16]);
  assign t[153] = (x[20] & x[21]);
  assign t[154] = (x[25] & x[26]);
  assign t[155] = (x[20] & x[30]);
  assign t[156] = (x[20] & x[32]);
  assign t[157] = (x[34] & x[35]);
  assign t[158] = (x[37] & x[38]);
  assign t[159] = (x[42] & x[43]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[160] = (x[25] & x[47]);
  assign t[161] = (x[25] & x[49]);
  assign t[162] = (x[51] & x[52]);
  assign t[163] = (x[56] & x[57]);
  assign t[164] = (x[20] & x[61]);
  assign t[165] = (x[34] & x[63]);
  assign t[166] = (x[34] & x[65]);
  assign t[167] = (x[37] & x[67]);
  assign t[168] = (x[37] & x[69]);
  assign t[169] = (x[42] & x[71]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (x[42] & x[73]);
  assign t[171] = (x[25] & x[75]);
  assign t[172] = (x[51] & x[77]);
  assign t[173] = (x[51] & x[79]);
  assign t[174] = (x[81] & x[82]);
  assign t[175] = (x[56] & x[84]);
  assign t[176] = (x[56] & x[86]);
  assign t[177] = (x[88] & x[89]);
  assign t[178] = (x[34] & x[91]);
  assign t[179] = (x[37] & x[93]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[180] = (x[42] & x[95]);
  assign t[181] = (x[51] & x[97]);
  assign t[182] = (x[81] & x[99]);
  assign t[183] = (x[81] & x[101]);
  assign t[184] = (x[56] & x[103]);
  assign t[185] = (x[88] & x[105]);
  assign t[186] = (x[88] & x[107]);
  assign t[187] = (x[81] & x[109]);
  assign t[188] = (x[88] & x[111]);
  assign t[18] = t[27] ^ t[28];
  assign t[19] = x[4] ? t[30] : t[29];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = t[35] ^ t[21];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[40] & t[41]);
  assign t[26] = ~(t[42] & t[112]);
  assign t[27] = t[43] ? x[24] : x[23];
  assign t[28] = ~(t[44] & t[45]);
  assign t[29] = ~(t[46] & t[47]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[48] ^ t[36];
  assign t[31] = ~(t[49] & t[50]);
  assign t[32] = t[51] ^ t[29];
  assign t[33] = ~(t[52] & t[53]);
  assign t[34] = ~(t[54] & t[113]);
  assign t[35] = t[110] ? x[29] : x[28];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[58];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[114]);
  assign t[41] = ~(t[115]);
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = ~(t[65]);
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = ~(t[68] & t[116]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[71] & t[117]);
  assign t[48] = t[43] ? x[41] : x[40];
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[74] & t[118]);
  assign t[51] = t[110] ? x[46] : x[45];
  assign t[52] = ~(t[119]);
  assign t[53] = ~(t[120]);
  assign t[54] = ~(t[75] & t[76]);
  assign t[55] = ~(t[77] & t[78]);
  assign t[56] = ~(t[79] & t[121]);
  assign t[57] = t[110] ? x[55] : x[54];
  assign t[58] = ~(t[80] & t[81]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[84] & t[122]);
  assign t[61] = t[43] ? x[60] : x[59];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = ~(t[115] & t[114]);
  assign t[64] = ~(t[123]);
  assign t[65] = ~(t[110]);
  assign t[66] = ~(t[124]);
  assign t[67] = ~(t[125]);
  assign t[68] = ~(t[87] & t[88]);
  assign t[69] = ~(t[126]);
  assign t[6] = ~(t[108] & t[109]);
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[89] & t[90]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[91] & t[92]);
  assign t[75] = ~(t[120] & t[119]);
  assign t[76] = ~(t[130]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[93] & t[94]);
  assign t[7] = ~(t[110] & t[111]);
  assign t[80] = ~(t[95] & t[96]);
  assign t[81] = ~(t[97] & t[133]);
  assign t[82] = ~(t[134]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[98] & t[99]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[136]);
  assign t[87] = ~(t[125] & t[124]);
  assign t[88] = ~(t[137]);
  assign t[89] = ~(t[127] & t[126]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[138]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[139]);
  assign t[93] = ~(t[132] & t[131]);
  assign t[94] = ~(t[140]);
  assign t[95] = ~(t[141]);
  assign t[96] = ~(t[142]);
  assign t[97] = ~(t[103] & t[104]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[143]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[107];
endmodule

module R1ind180(x, y);
 input [94:0] x;
 output y;

 wire [154:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[132] ^ x[35];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[40];
  assign t[103] = t[135] ^ x[43];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[50];
  assign t[106] = t[138] ^ x[52];
  assign t[107] = t[139] ^ x[56];
  assign t[108] = t[140] ^ x[59];
  assign t[109] = t[141] ^ x[61];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[142] ^ x[66];
  assign t[111] = t[143] ^ x[68];
  assign t[112] = t[144] ^ x[72];
  assign t[113] = t[145] ^ x[74];
  assign t[114] = t[146] ^ x[76];
  assign t[115] = t[147] ^ x[78];
  assign t[116] = t[148] ^ x[81];
  assign t[117] = t[149] ^ x[83];
  assign t[118] = t[150] ^ x[85];
  assign t[119] = t[151] ^ x[88];
  assign t[11] = t[94] ? x[18] : x[19];
  assign t[120] = t[152] ^ x[90];
  assign t[121] = t[153] ^ x[92];
  assign t[122] = t[154] ^ x[94];
  assign t[123] = (x[0] & x[1]);
  assign t[124] = (x[6] & x[7]);
  assign t[125] = (x[9] & x[10]);
  assign t[126] = (x[12] & x[13]);
  assign t[127] = (x[15] & x[16]);
  assign t[128] = (x[20] & x[21]);
  assign t[129] = (x[20] & x[23]);
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = (x[27] & x[28]);
  assign t[131] = (x[27] & x[30]);
  assign t[132] = (x[20] & x[34]);
  assign t[133] = (x[36] & x[37]);
  assign t[134] = (x[36] & x[39]);
  assign t[135] = (x[41] & x[42]);
  assign t[136] = (x[41] & x[44]);
  assign t[137] = (x[48] & x[49]);
  assign t[138] = (x[48] & x[51]);
  assign t[139] = (x[27] & x[55]);
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (x[57] & x[58]);
  assign t[141] = (x[57] & x[60]);
  assign t[142] = (x[64] & x[65]);
  assign t[143] = (x[64] & x[67]);
  assign t[144] = (x[36] & x[71]);
  assign t[145] = (x[41] & x[73]);
  assign t[146] = (x[48] & x[75]);
  assign t[147] = (x[57] & x[77]);
  assign t[148] = (x[79] & x[80]);
  assign t[149] = (x[79] & x[82]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[64] & x[84]);
  assign t[151] = (x[86] & x[87]);
  assign t[152] = (x[86] & x[89]);
  assign t[153] = (x[79] & x[91]);
  assign t[154] = (x[86] & x[93]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = t[27] ^ t[28];
  assign t[19] = x[4] ? t[30] : t[29];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = t[35] ^ t[21];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[96] & t[40]);
  assign t[26] = ~(t[97] & t[41]);
  assign t[27] = t[42] ? x[26] : x[25];
  assign t[28] = ~(t[43] & t[44]);
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[47] ^ t[31];
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[36];
  assign t[33] = ~(t[98] & t[51]);
  assign t[34] = ~(t[99] & t[52]);
  assign t[35] = t[94] ? x[33] : x[32];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = t[55] ^ t[56];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[100]);
  assign t[41] = ~(t[100] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[101] & t[63]);
  assign t[44] = ~(t[102] & t[64]);
  assign t[45] = ~(t[103] & t[65]);
  assign t[46] = ~(t[104] & t[66]);
  assign t[47] = t[67] ? x[47] : x[46];
  assign t[48] = ~(t[105] & t[68]);
  assign t[49] = ~(t[106] & t[69]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[70] ? x[54] : x[53];
  assign t[51] = ~(t[107]);
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = ~(t[109] & t[73]);
  assign t[55] = t[94] ? x[63] : x[62];
  assign t[56] = ~(t[74] & t[75]);
  assign t[57] = ~(t[110] & t[76]);
  assign t[58] = ~(t[111] & t[77]);
  assign t[59] = t[42] ? x[70] : x[69];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[78] & t[79]);
  assign t[61] = ~(t[96]);
  assign t[62] = ~(t[94]);
  assign t[63] = ~(t[112]);
  assign t[64] = ~(t[112] & t[80]);
  assign t[65] = ~(t[113]);
  assign t[66] = ~(t[113] & t[81]);
  assign t[67] = ~(t[62]);
  assign t[68] = ~(t[114]);
  assign t[69] = ~(t[114] & t[82]);
  assign t[6] = ~(t[92] & t[93]);
  assign t[70] = ~(t[62]);
  assign t[71] = ~(t[98]);
  assign t[72] = ~(t[115]);
  assign t[73] = ~(t[115] & t[83]);
  assign t[74] = ~(t[116] & t[84]);
  assign t[75] = ~(t[117] & t[85]);
  assign t[76] = ~(t[118]);
  assign t[77] = ~(t[118] & t[86]);
  assign t[78] = ~(t[119] & t[87]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[94] & t[95]);
  assign t[80] = ~(t[101]);
  assign t[81] = ~(t[103]);
  assign t[82] = ~(t[105]);
  assign t[83] = ~(t[108]);
  assign t[84] = ~(t[121]);
  assign t[85] = ~(t[121] & t[89]);
  assign t[86] = ~(t[110]);
  assign t[87] = ~(t[122]);
  assign t[88] = ~(t[122] & t[90]);
  assign t[89] = ~(t[116]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[119]);
  assign t[91] = t[123] ^ x[2];
  assign t[92] = t[124] ^ x[8];
  assign t[93] = t[125] ^ x[11];
  assign t[94] = t[126] ^ x[14];
  assign t[95] = t[127] ^ x[17];
  assign t[96] = t[128] ^ x[22];
  assign t[97] = t[129] ^ x[24];
  assign t[98] = t[130] ^ x[29];
  assign t[99] = t[131] ^ x[31];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[91];
endmodule

module R1ind181(x, y);
 input [112:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[212] | t[213]);
  assign t[101] = ~(t[137] & t[139]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[140] | t[141]);
  assign t[105] = ~(t[142] | t[143]);
  assign t[106] = ~(t[226] | t[144]);
  assign t[107] = t[203] ? x[81] : x[80];
  assign t[108] = ~(t[145] & t[146]);
  assign t[109] = ~(t[227]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = ~(t[228]);
  assign t[111] = ~(t[147] | t[148]);
  assign t[112] = ~(t[149] | t[150]);
  assign t[113] = ~(t[229] | t[151]);
  assign t[114] = t[203] ? x[90] : x[89];
  assign t[115] = ~(t[145] & t[152]);
  assign t[116] = ~(t[121] | t[201]);
  assign t[117] = ~(t[153] & t[154]);
  assign t[118] = ~(t[202] | t[155]);
  assign t[119] = t[79] & t[201];
  assign t[11] = ~(t[15] ^ t[16]);
  assign t[120] = ~(t[121] | t[156]);
  assign t[121] = ~(t[203]);
  assign t[122] = t[201] ? t[158] : t[157];
  assign t[123] = ~(t[159] & t[204]);
  assign t[124] = ~(t[160] & t[155]);
  assign t[125] = ~(t[230]);
  assign t[126] = ~(t[217] | t[218]);
  assign t[127] = ~(t[161] & t[162]);
  assign t[128] = ~(t[163] & t[78]);
  assign t[129] = ~(t[79] | t[164]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[130] = ~(t[79] | t[165]);
  assign t[131] = ~(t[231]);
  assign t[132] = ~(t[219] | t[220]);
  assign t[133] = ~(t[129] | t[166]);
  assign t[134] = ~(t[167] | t[168]);
  assign t[135] = ~(t[232]);
  assign t[136] = ~(t[221] | t[222]);
  assign t[137] = ~(t[48] | t[169]);
  assign t[138] = ~(t[170] | t[171]);
  assign t[139] = ~(t[166] | t[130]);
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = ~(t[233]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[234]);
  assign t[143] = ~(t[235]);
  assign t[144] = ~(t[172] | t[173]);
  assign t[145] = ~(t[48] | t[174]);
  assign t[146] = ~(t[120] | t[175]);
  assign t[147] = ~(t[236]);
  assign t[148] = ~(t[227] | t[228]);
  assign t[149] = ~(t[237]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = ~(t[238]);
  assign t[151] = ~(t[176] | t[177]);
  assign t[152] = ~(t[178] | t[130]);
  assign t[153] = ~(t[204] & t[179]);
  assign t[154] = ~(x[4] & t[118]);
  assign t[155] = ~(t[204]);
  assign t[156] = t[201] ? t[157] : t[158];
  assign t[157] = ~(t[179] & t[155]);
  assign t[158] = ~(x[4] & t[180]);
  assign t[159] = x[4] & t[202];
  assign t[15] = x[4] ? t[24] : t[23];
  assign t[160] = ~(x[4] | t[202]);
  assign t[161] = ~(t[170] | t[181]);
  assign t[162] = ~(t[121] & t[182]);
  assign t[163] = ~(t[183] & t[184]);
  assign t[164] = t[201] ? t[123] : t[124];
  assign t[165] = t[201] ? t[186] : t[185];
  assign t[166] = ~(t[79] | t[187]);
  assign t[167] = t[171] | t[188];
  assign t[168] = ~(t[189] & t[78]);
  assign t[169] = ~(t[79] | t[190]);
  assign t[16] = ~(t[25] ^ t[26]);
  assign t[170] = ~(t[121] | t[191]);
  assign t[171] = ~(t[192] & t[76]);
  assign t[172] = ~(t[239]);
  assign t[173] = ~(t[234] | t[235]);
  assign t[174] = ~(t[133] & t[163]);
  assign t[175] = t[169] | t[193];
  assign t[176] = ~(t[240]);
  assign t[177] = ~(t[237] | t[238]);
  assign t[178] = ~(t[79] | t[194]);
  assign t[179] = ~(x[4] | t[195]);
  assign t[17] = t[27] ? x[18] : x[19];
  assign t[180] = ~(t[202] | t[204]);
  assign t[181] = ~(t[79] | t[196]);
  assign t[182] = ~(t[158] & t[153]);
  assign t[183] = t[204] & t[116];
  assign t[184] = t[160] | t[159];
  assign t[185] = ~(t[160] & t[204]);
  assign t[186] = ~(t[159] & t[155]);
  assign t[187] = t[201] ? t[158] : t[153];
  assign t[188] = ~(t[79] | t[197]);
  assign t[189] = ~(t[193] | t[178]);
  assign t[18] = ~(t[28] & t[29]);
  assign t[190] = t[201] ? t[185] : t[186];
  assign t[191] = t[201] ? t[124] : t[186];
  assign t[192] = ~(t[198] | t[120]);
  assign t[193] = ~(t[75]);
  assign t[194] = t[201] ? t[154] : t[157];
  assign t[195] = ~(t[202]);
  assign t[196] = t[201] ? t[157] : t[154];
  assign t[197] = t[201] ? t[153] : t[158];
  assign t[198] = ~(t[121] | t[199]);
  assign t[199] = t[201] ? t[186] : t[124];
  assign t[19] = ~(t[30] | t[31]);
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[200] = t[241] ^ x[2];
  assign t[201] = t[242] ^ x[8];
  assign t[202] = t[243] ^ x[11];
  assign t[203] = t[244] ^ x[14];
  assign t[204] = t[245] ^ x[17];
  assign t[205] = t[246] ^ x[22];
  assign t[206] = t[247] ^ x[25];
  assign t[207] = t[248] ^ x[27];
  assign t[208] = t[249] ^ x[29];
  assign t[209] = t[250] ^ x[32];
  assign t[20] = ~(t[32] ^ t[33]);
  assign t[210] = t[251] ^ x[37];
  assign t[211] = t[252] ^ x[40];
  assign t[212] = t[253] ^ x[42];
  assign t[213] = t[254] ^ x[44];
  assign t[214] = t[255] ^ x[49];
  assign t[215] = t[256] ^ x[52];
  assign t[216] = t[257] ^ x[54];
  assign t[217] = t[258] ^ x[56];
  assign t[218] = t[259] ^ x[58];
  assign t[219] = t[260] ^ x[60];
  assign t[21] = x[4] ? t[35] : t[34];
  assign t[220] = t[261] ^ x[62];
  assign t[221] = t[262] ^ x[66];
  assign t[222] = t[263] ^ x[68];
  assign t[223] = t[264] ^ x[72];
  assign t[224] = t[265] ^ x[74];
  assign t[225] = t[266] ^ x[76];
  assign t[226] = t[267] ^ x[79];
  assign t[227] = t[268] ^ x[83];
  assign t[228] = t[269] ^ x[85];
  assign t[229] = t[270] ^ x[88];
  assign t[22] = x[4] ? t[37] : t[36];
  assign t[230] = t[271] ^ x[92];
  assign t[231] = t[272] ^ x[94];
  assign t[232] = t[273] ^ x[96];
  assign t[233] = t[274] ^ x[98];
  assign t[234] = t[275] ^ x[100];
  assign t[235] = t[276] ^ x[102];
  assign t[236] = t[277] ^ x[104];
  assign t[237] = t[278] ^ x[106];
  assign t[238] = t[279] ^ x[108];
  assign t[239] = t[280] ^ x[110];
  assign t[23] = ~(t[38] | t[39]);
  assign t[240] = t[281] ^ x[112];
  assign t[241] = (x[0] & x[1]);
  assign t[242] = (x[6] & x[7]);
  assign t[243] = (x[9] & x[10]);
  assign t[244] = (x[12] & x[13]);
  assign t[245] = (x[15] & x[16]);
  assign t[246] = (x[20] & x[21]);
  assign t[247] = (x[23] & x[24]);
  assign t[248] = (x[20] & x[26]);
  assign t[249] = (x[20] & x[28]);
  assign t[24] = ~(t[23] ^ t[40]);
  assign t[250] = (x[30] & x[31]);
  assign t[251] = (x[35] & x[36]);
  assign t[252] = (x[38] & x[39]);
  assign t[253] = (x[23] & x[41]);
  assign t[254] = (x[23] & x[43]);
  assign t[255] = (x[47] & x[48]);
  assign t[256] = (x[50] & x[51]);
  assign t[257] = (x[20] & x[53]);
  assign t[258] = (x[30] & x[55]);
  assign t[259] = (x[30] & x[57]);
  assign t[25] = x[4] ? t[42] : t[41];
  assign t[260] = (x[35] & x[59]);
  assign t[261] = (x[35] & x[61]);
  assign t[262] = (x[38] & x[65]);
  assign t[263] = (x[38] & x[67]);
  assign t[264] = (x[23] & x[71]);
  assign t[265] = (x[47] & x[73]);
  assign t[266] = (x[47] & x[75]);
  assign t[267] = (x[77] & x[78]);
  assign t[268] = (x[50] & x[82]);
  assign t[269] = (x[50] & x[84]);
  assign t[26] = x[4] ? t[44] : t[43];
  assign t[270] = (x[86] & x[87]);
  assign t[271] = (x[30] & x[91]);
  assign t[272] = (x[35] & x[93]);
  assign t[273] = (x[38] & x[95]);
  assign t[274] = (x[47] & x[97]);
  assign t[275] = (x[77] & x[99]);
  assign t[276] = (x[77] & x[101]);
  assign t[277] = (x[50] & x[103]);
  assign t[278] = (x[86] & x[105]);
  assign t[279] = (x[86] & x[107]);
  assign t[27] = ~(t[45]);
  assign t[280] = (x[77] & x[109]);
  assign t[281] = (x[86] & x[111]);
  assign t[28] = ~(t[46] | t[47]);
  assign t[29] = ~(t[48]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[205] | t[51]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[33] = ~(t[54] ^ t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[43] ^ t[58]);
  assign t[36] = ~(t[59] | t[60]);
  assign t[37] = ~(t[34] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[206] | t[64]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[65] ^ t[66]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[42] = ~(t[69] ^ t[70]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[45] = ~(t[203]);
  assign t[46] = ~(t[75] & t[76]);
  assign t[47] = ~(t[77] & t[78]);
  assign t[48] = ~(t[79] | t[80]);
  assign t[49] = ~(t[207]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[208]);
  assign t[51] = ~(t[81] | t[82]);
  assign t[52] = ~(t[83] | t[84]);
  assign t[53] = ~(t[209] | t[85]);
  assign t[54] = t[86] ? x[34] : x[33];
  assign t[55] = ~(t[87] & t[88]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[210] | t[91]);
  assign t[58] = ~(t[92] ^ t[93]);
  assign t[59] = ~(t[94] | t[95]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[211] | t[96]);
  assign t[61] = ~(t[97] ^ t[98]);
  assign t[62] = ~(t[212]);
  assign t[63] = ~(t[213]);
  assign t[64] = ~(t[99] | t[100]);
  assign t[65] = t[203] ? x[46] : x[45];
  assign t[66] = t[46] | t[101];
  assign t[67] = ~(t[102] | t[103]);
  assign t[68] = ~(t[214] | t[104]);
  assign t[69] = ~(t[105] | t[106]);
  assign t[6] = ~(t[201] & t[202]);
  assign t[70] = ~(t[107] ^ t[108]);
  assign t[71] = ~(t[109] | t[110]);
  assign t[72] = ~(t[215] | t[111]);
  assign t[73] = ~(t[112] | t[113]);
  assign t[74] = ~(t[114] ^ t[115]);
  assign t[75] = ~(t[116] & t[117]);
  assign t[76] = ~(t[118] & t[119]);
  assign t[77] = ~(t[120]);
  assign t[78] = t[121] | t[122];
  assign t[79] = ~(t[121]);
  assign t[7] = ~(t[203] & t[204]);
  assign t[80] = t[201] ? t[124] : t[123];
  assign t[81] = ~(t[216]);
  assign t[82] = ~(t[207] | t[208]);
  assign t[83] = ~(t[217]);
  assign t[84] = ~(t[218]);
  assign t[85] = ~(t[125] | t[126]);
  assign t[86] = ~(t[45]);
  assign t[87] = ~(t[127] | t[128]);
  assign t[88] = ~(t[129] | t[130]);
  assign t[89] = ~(t[219]);
  assign t[8] = ~(t[11] ^ t[12]);
  assign t[90] = ~(t[220]);
  assign t[91] = ~(t[131] | t[132]);
  assign t[92] = t[86] ? x[64] : x[63];
  assign t[93] = ~(t[133] & t[134]);
  assign t[94] = ~(t[221]);
  assign t[95] = ~(t[222]);
  assign t[96] = ~(t[135] | t[136]);
  assign t[97] = t[86] ? x[70] : x[69];
  assign t[98] = ~(t[137] & t[138]);
  assign t[99] = ~(t[223]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[200];
endmodule

module R1ind182(x, y);
 input [79:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = (x[20] & x[21]);
  assign t[101] = (x[20] & x[25]);
  assign t[102] = (x[20] & x[27]);
  assign t[103] = (x[29] & x[30]);
  assign t[104] = (x[32] & x[33]);
  assign t[105] = (x[37] & x[38]);
  assign t[106] = (x[20] & x[42]);
  assign t[107] = (x[29] & x[44]);
  assign t[108] = (x[29] & x[46]);
  assign t[109] = (x[32] & x[48]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = (x[32] & x[50]);
  assign t[111] = (x[52] & x[53]);
  assign t[112] = (x[37] & x[55]);
  assign t[113] = (x[37] & x[57]);
  assign t[114] = (x[59] & x[60]);
  assign t[115] = (x[29] & x[62]);
  assign t[116] = (x[32] & x[64]);
  assign t[117] = (x[52] & x[66]);
  assign t[118] = (x[52] & x[68]);
  assign t[119] = (x[37] & x[70]);
  assign t[11] = t[69] ? x[18] : x[19];
  assign t[120] = (x[59] & x[72]);
  assign t[121] = (x[59] & x[74]);
  assign t[122] = (x[52] & x[76]);
  assign t[123] = (x[59] & x[78]);
  assign t[12] = x[4] ? t[15] : t[14];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = t[20] ^ t[21];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = t[28] | t[71];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[69] ? x[24] : x[23];
  assign t[21] = ~(t[29] & t[30]);
  assign t[22] = ~(t[31] & t[32]);
  assign t[23] = t[33] ^ t[34];
  assign t[24] = ~(t[35] & t[36]);
  assign t[25] = t[37] ^ t[38];
  assign t[26] = ~(t[72]);
  assign t[27] = ~(t[73]);
  assign t[28] = ~(t[39] | t[26]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[42] | t[74];
  assign t[31] = ~(t[43] & t[44]);
  assign t[32] = t[45] | t[75];
  assign t[33] = t[69] ? x[36] : x[35];
  assign t[34] = ~(t[46] & t[47]);
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = t[50] | t[76];
  assign t[37] = t[51] ? x[41] : x[40];
  assign t[38] = ~(t[52] & t[53]);
  assign t[39] = ~(t[77]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[78]);
  assign t[41] = ~(t[79]);
  assign t[42] = ~(t[54] | t[40]);
  assign t[43] = ~(t[80]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[55] | t[43]);
  assign t[46] = ~(t[56] & t[57]);
  assign t[47] = t[58] | t[82];
  assign t[48] = ~(t[83]);
  assign t[49] = ~(t[84]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[59] | t[48]);
  assign t[51] = ~(t[60]);
  assign t[52] = ~(t[61] & t[62]);
  assign t[53] = t[63] | t[85];
  assign t[54] = ~(t[86]);
  assign t[55] = ~(t[87]);
  assign t[56] = ~(t[88]);
  assign t[57] = ~(t[89]);
  assign t[58] = ~(t[64] | t[56]);
  assign t[59] = ~(t[90]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[69]);
  assign t[61] = ~(t[91]);
  assign t[62] = ~(t[92]);
  assign t[63] = ~(t[65] | t[61]);
  assign t[64] = ~(t[93]);
  assign t[65] = ~(t[94]);
  assign t[66] = t[95] ^ x[2];
  assign t[67] = t[96] ^ x[8];
  assign t[68] = t[97] ^ x[11];
  assign t[69] = t[98] ^ x[14];
  assign t[6] = ~(t[67] & t[68]);
  assign t[70] = t[99] ^ x[17];
  assign t[71] = t[100] ^ x[22];
  assign t[72] = t[101] ^ x[26];
  assign t[73] = t[102] ^ x[28];
  assign t[74] = t[103] ^ x[31];
  assign t[75] = t[104] ^ x[34];
  assign t[76] = t[105] ^ x[39];
  assign t[77] = t[106] ^ x[43];
  assign t[78] = t[107] ^ x[45];
  assign t[79] = t[108] ^ x[47];
  assign t[7] = ~(t[69] & t[70]);
  assign t[80] = t[109] ^ x[49];
  assign t[81] = t[110] ^ x[51];
  assign t[82] = t[111] ^ x[54];
  assign t[83] = t[112] ^ x[56];
  assign t[84] = t[113] ^ x[58];
  assign t[85] = t[114] ^ x[61];
  assign t[86] = t[115] ^ x[63];
  assign t[87] = t[116] ^ x[65];
  assign t[88] = t[117] ^ x[67];
  assign t[89] = t[118] ^ x[69];
  assign t[8] = t[11] ^ t[9];
  assign t[90] = t[119] ^ x[71];
  assign t[91] = t[120] ^ x[73];
  assign t[92] = t[121] ^ x[75];
  assign t[93] = t[122] ^ x[77];
  assign t[94] = t[123] ^ x[79];
  assign t[95] = (x[0] & x[1]);
  assign t[96] = (x[6] & x[7]);
  assign t[97] = (x[9] & x[10]);
  assign t[98] = (x[12] & x[13]);
  assign t[99] = (x[15] & x[16]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = t[0] ? t[1] : t[66];
endmodule

module R1ind183(x, y);
 input [79:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[129] ^ x[79];
  assign t[101] = (x[0] & x[1]);
  assign t[102] = (x[6] & x[7]);
  assign t[103] = (x[9] & x[10]);
  assign t[104] = (x[12] & x[13]);
  assign t[105] = (x[15] & x[16]);
  assign t[106] = (x[20] & x[21]);
  assign t[107] = (x[20] & x[25]);
  assign t[108] = (x[20] & x[27]);
  assign t[109] = (x[29] & x[30]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = (x[32] & x[33]);
  assign t[111] = (x[37] & x[38]);
  assign t[112] = (x[20] & x[42]);
  assign t[113] = (x[29] & x[44]);
  assign t[114] = (x[29] & x[46]);
  assign t[115] = (x[32] & x[48]);
  assign t[116] = (x[32] & x[50]);
  assign t[117] = (x[52] & x[53]);
  assign t[118] = (x[37] & x[55]);
  assign t[119] = (x[37] & x[57]);
  assign t[11] = t[75] ? x[18] : x[19];
  assign t[120] = (x[59] & x[60]);
  assign t[121] = (x[29] & x[62]);
  assign t[122] = (x[32] & x[64]);
  assign t[123] = (x[52] & x[66]);
  assign t[124] = (x[52] & x[68]);
  assign t[125] = (x[37] & x[70]);
  assign t[126] = (x[59] & x[72]);
  assign t[127] = (x[59] & x[74]);
  assign t[128] = (x[52] & x[76]);
  assign t[129] = (x[59] & x[78]);
  assign t[12] = x[4] ? t[15] : t[14];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = t[20] ^ t[21];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[77]);
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[75] ? x[24] : x[23];
  assign t[21] = ~(t[29] & t[30]);
  assign t[22] = ~(t[31] & t[32]);
  assign t[23] = t[33] ^ t[34];
  assign t[24] = ~(t[35] & t[36]);
  assign t[25] = t[37] ^ t[38];
  assign t[26] = ~(t[78]);
  assign t[27] = ~(t[79]);
  assign t[28] = ~(t[39] & t[40]);
  assign t[29] = ~(t[41] & t[42]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[43] & t[80]);
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = ~(t[46] & t[81]);
  assign t[33] = t[75] ? x[36] : x[35];
  assign t[34] = ~(t[47] & t[48]);
  assign t[35] = ~(t[49] & t[50]);
  assign t[36] = ~(t[51] & t[82]);
  assign t[37] = t[52] ? x[41] : x[40];
  assign t[38] = ~(t[53] & t[54]);
  assign t[39] = ~(t[79] & t[78]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[83]);
  assign t[41] = ~(t[84]);
  assign t[42] = ~(t[85]);
  assign t[43] = ~(t[55] & t[56]);
  assign t[44] = ~(t[86]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[57] & t[58]);
  assign t[47] = ~(t[59] & t[60]);
  assign t[48] = ~(t[61] & t[88]);
  assign t[49] = ~(t[89]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[90]);
  assign t[51] = ~(t[62] & t[63]);
  assign t[52] = ~(t[64]);
  assign t[53] = ~(t[65] & t[66]);
  assign t[54] = ~(t[67] & t[91]);
  assign t[55] = ~(t[85] & t[84]);
  assign t[56] = ~(t[92]);
  assign t[57] = ~(t[87] & t[86]);
  assign t[58] = ~(t[93]);
  assign t[59] = ~(t[94]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[95]);
  assign t[61] = ~(t[68] & t[69]);
  assign t[62] = ~(t[90] & t[89]);
  assign t[63] = ~(t[96]);
  assign t[64] = ~(t[75]);
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[70] & t[71]);
  assign t[68] = ~(t[95] & t[94]);
  assign t[69] = ~(t[99]);
  assign t[6] = ~(t[73] & t[74]);
  assign t[70] = ~(t[98] & t[97]);
  assign t[71] = ~(t[100]);
  assign t[72] = t[101] ^ x[2];
  assign t[73] = t[102] ^ x[8];
  assign t[74] = t[103] ^ x[11];
  assign t[75] = t[104] ^ x[14];
  assign t[76] = t[105] ^ x[17];
  assign t[77] = t[106] ^ x[22];
  assign t[78] = t[107] ^ x[26];
  assign t[79] = t[108] ^ x[28];
  assign t[7] = ~(t[75] & t[76]);
  assign t[80] = t[109] ^ x[31];
  assign t[81] = t[110] ^ x[34];
  assign t[82] = t[111] ^ x[39];
  assign t[83] = t[112] ^ x[43];
  assign t[84] = t[113] ^ x[45];
  assign t[85] = t[114] ^ x[47];
  assign t[86] = t[115] ^ x[49];
  assign t[87] = t[116] ^ x[51];
  assign t[88] = t[117] ^ x[54];
  assign t[89] = t[118] ^ x[56];
  assign t[8] = t[11] ^ t[9];
  assign t[90] = t[119] ^ x[58];
  assign t[91] = t[120] ^ x[61];
  assign t[92] = t[121] ^ x[63];
  assign t[93] = t[122] ^ x[65];
  assign t[94] = t[123] ^ x[67];
  assign t[95] = t[124] ^ x[69];
  assign t[96] = t[125] ^ x[71];
  assign t[97] = t[126] ^ x[73];
  assign t[98] = t[127] ^ x[75];
  assign t[99] = t[128] ^ x[77];
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = t[0] ? t[1] : t[72];
endmodule

module R1ind184(x, y);
 input [67:0] x;
 output y;

 wire [105:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = (x[52] & x[55]);
  assign t[101] = (x[41] & x[57]);
  assign t[102] = (x[59] & x[60]);
  assign t[103] = (x[59] & x[62]);
  assign t[104] = (x[52] & x[64]);
  assign t[105] = (x[59] & x[66]);
  assign t[10] = x[18] ^ x[19];
  assign t[11] = t[63] ? x[19] : x[18];
  assign t[12] = x[4] ? t[15] : t[14];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[14] = ~(t[18] & t[19]);
  assign t[15] = t[20] ^ t[21];
  assign t[16] = x[4] ? t[23] : t[22];
  assign t[17] = x[4] ? t[25] : t[24];
  assign t[18] = ~(t[65] & t[26]);
  assign t[19] = ~(t[66] & t[27]);
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[63] ? x[26] : x[25];
  assign t[21] = ~(t[28] & t[29]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = t[32] ^ t[33];
  assign t[24] = ~(t[34] & t[35]);
  assign t[25] = t[36] ^ t[37];
  assign t[26] = ~(t[67]);
  assign t[27] = ~(t[67] & t[38]);
  assign t[28] = ~(t[68] & t[39]);
  assign t[29] = ~(t[69] & t[40]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[70] & t[41]);
  assign t[31] = ~(t[71] & t[42]);
  assign t[32] = t[63] ? x[40] : x[39];
  assign t[33] = ~(t[43] & t[44]);
  assign t[34] = ~(t[72] & t[45]);
  assign t[35] = ~(t[73] & t[46]);
  assign t[36] = t[47] ? x[47] : x[46];
  assign t[37] = ~(t[48] & t[49]);
  assign t[38] = ~(t[65]);
  assign t[39] = ~(t[74]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[74] & t[50]);
  assign t[41] = ~(t[75]);
  assign t[42] = ~(t[75] & t[51]);
  assign t[43] = ~(t[76] & t[52]);
  assign t[44] = ~(t[77] & t[53]);
  assign t[45] = ~(t[78]);
  assign t[46] = ~(t[78] & t[54]);
  assign t[47] = ~(t[55]);
  assign t[48] = ~(t[79] & t[56]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[68]);
  assign t[51] = ~(t[70]);
  assign t[52] = ~(t[81]);
  assign t[53] = ~(t[81] & t[58]);
  assign t[54] = ~(t[72]);
  assign t[55] = ~(t[63]);
  assign t[56] = ~(t[82]);
  assign t[57] = ~(t[82] & t[59]);
  assign t[58] = ~(t[76]);
  assign t[59] = ~(t[79]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = t[83] ^ x[2];
  assign t[61] = t[84] ^ x[8];
  assign t[62] = t[85] ^ x[11];
  assign t[63] = t[86] ^ x[14];
  assign t[64] = t[87] ^ x[17];
  assign t[65] = t[88] ^ x[22];
  assign t[66] = t[89] ^ x[24];
  assign t[67] = t[90] ^ x[28];
  assign t[68] = t[91] ^ x[31];
  assign t[69] = t[92] ^ x[33];
  assign t[6] = ~(t[61] & t[62]);
  assign t[70] = t[93] ^ x[36];
  assign t[71] = t[94] ^ x[38];
  assign t[72] = t[95] ^ x[43];
  assign t[73] = t[96] ^ x[45];
  assign t[74] = t[97] ^ x[49];
  assign t[75] = t[98] ^ x[51];
  assign t[76] = t[99] ^ x[54];
  assign t[77] = t[100] ^ x[56];
  assign t[78] = t[101] ^ x[58];
  assign t[79] = t[102] ^ x[61];
  assign t[7] = ~(t[63] & t[64]);
  assign t[80] = t[103] ^ x[63];
  assign t[81] = t[104] ^ x[65];
  assign t[82] = t[105] ^ x[67];
  assign t[83] = (x[0] & x[1]);
  assign t[84] = (x[6] & x[7]);
  assign t[85] = (x[9] & x[10]);
  assign t[86] = (x[12] & x[13]);
  assign t[87] = (x[15] & x[16]);
  assign t[88] = (x[20] & x[21]);
  assign t[89] = (x[20] & x[23]);
  assign t[8] = t[11] ^ t[9];
  assign t[90] = (x[20] & x[27]);
  assign t[91] = (x[29] & x[30]);
  assign t[92] = (x[29] & x[32]);
  assign t[93] = (x[34] & x[35]);
  assign t[94] = (x[34] & x[37]);
  assign t[95] = (x[41] & x[42]);
  assign t[96] = (x[41] & x[44]);
  assign t[97] = (x[29] & x[48]);
  assign t[98] = (x[34] & x[50]);
  assign t[99] = (x[52] & x[53]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = t[0] ? t[1] : t[60];
endmodule

module R1ind185(x, y);
 input [79:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[153] | t[154]);
  assign t[101] = ~(t[161]);
  assign t[102] = ~(t[162]);
  assign t[103] = ~(t[118] | t[119]);
  assign t[104] = ~(t[120] | t[56]);
  assign t[105] = ~(x[4] | t[121]);
  assign t[106] = ~(t[122] & t[140]);
  assign t[107] = ~(t[123] & t[82]);
  assign t[108] = ~(t[122] & t[82]);
  assign t[109] = ~(t[123] & t[140]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = ~(x[4] & t[124]);
  assign t[111] = ~(t[116]);
  assign t[112] = t[79] | t[125];
  assign t[113] = ~(t[163]);
  assign t[114] = ~(t[158] | t[159]);
  assign t[115] = ~(t[126] & t[127]);
  assign t[116] = ~(t[79] | t[128]);
  assign t[117] = t[54] | t[129];
  assign t[118] = ~(t[164]);
  assign t[119] = ~(t[161] | t[162]);
  assign t[11] = ~(t[14] ^ t[15]);
  assign t[120] = ~(t[83] | t[130]);
  assign t[121] = ~(t[138]);
  assign t[122] = x[4] & t[138];
  assign t[123] = ~(x[4] | t[138]);
  assign t[124] = ~(t[138] | t[140]);
  assign t[125] = t[137] ? t[110] : t[131];
  assign t[126] = ~(t[132] | t[55]);
  assign t[127] = ~(t[133] & t[134]);
  assign t[128] = t[137] ? t[131] : t[110];
  assign t[129] = ~(t[30]);
  assign t[12] = x[4] ? t[17] : t[16];
  assign t[130] = t[137] ? t[81] : t[131];
  assign t[131] = ~(t[105] & t[82]);
  assign t[132] = ~(t[83] | t[135]);
  assign t[133] = t[140] & t[49];
  assign t[134] = t[123] | t[122];
  assign t[135] = t[137] ? t[106] : t[107];
  assign t[136] = t[165] ^ x[2];
  assign t[137] = t[166] ^ x[8];
  assign t[138] = t[167] ^ x[11];
  assign t[139] = t[168] ^ x[14];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[169] ^ x[17];
  assign t[141] = t[170] ^ x[22];
  assign t[142] = t[171] ^ x[24];
  assign t[143] = t[172] ^ x[26];
  assign t[144] = t[173] ^ x[29];
  assign t[145] = t[174] ^ x[34];
  assign t[146] = t[175] ^ x[37];
  assign t[147] = t[176] ^ x[39];
  assign t[148] = t[177] ^ x[41];
  assign t[149] = t[178] ^ x[43];
  assign t[14] = t[139] ? x[19] : x[18];
  assign t[150] = t[179] ^ x[45];
  assign t[151] = t[180] ^ x[47];
  assign t[152] = t[181] ^ x[50];
  assign t[153] = t[182] ^ x[54];
  assign t[154] = t[183] ^ x[56];
  assign t[155] = t[184] ^ x[59];
  assign t[156] = t[185] ^ x[63];
  assign t[157] = t[186] ^ x[65];
  assign t[158] = t[187] ^ x[67];
  assign t[159] = t[188] ^ x[69];
  assign t[15] = t[20] | t[21];
  assign t[160] = t[189] ^ x[71];
  assign t[161] = t[190] ^ x[73];
  assign t[162] = t[191] ^ x[75];
  assign t[163] = t[192] ^ x[77];
  assign t[164] = t[193] ^ x[79];
  assign t[165] = (x[0] & x[1]);
  assign t[166] = (x[6] & x[7]);
  assign t[167] = (x[9] & x[10]);
  assign t[168] = (x[12] & x[13]);
  assign t[169] = (x[15] & x[16]);
  assign t[16] = ~(t[22] | t[23]);
  assign t[170] = (x[20] & x[21]);
  assign t[171] = (x[20] & x[23]);
  assign t[172] = (x[20] & x[25]);
  assign t[173] = (x[27] & x[28]);
  assign t[174] = (x[32] & x[33]);
  assign t[175] = (x[35] & x[36]);
  assign t[176] = (x[20] & x[38]);
  assign t[177] = (x[27] & x[40]);
  assign t[178] = (x[27] & x[42]);
  assign t[179] = (x[32] & x[44]);
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = (x[32] & x[46]);
  assign t[181] = (x[48] & x[49]);
  assign t[182] = (x[35] & x[53]);
  assign t[183] = (x[35] & x[55]);
  assign t[184] = (x[57] & x[58]);
  assign t[185] = (x[27] & x[62]);
  assign t[186] = (x[32] & x[64]);
  assign t[187] = (x[48] & x[66]);
  assign t[188] = (x[48] & x[68]);
  assign t[189] = (x[35] & x[70]);
  assign t[18] = x[4] ? t[27] : t[26];
  assign t[190] = (x[57] & x[72]);
  assign t[191] = (x[57] & x[74]);
  assign t[192] = (x[48] & x[76]);
  assign t[193] = (x[57] & x[78]);
  assign t[19] = x[4] ? t[29] : t[28];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = ~(t[30] & t[31]);
  assign t[21] = ~(t[32] & t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[141] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = ~(t[39] ^ t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[28] = ~(t[45] | t[46]);
  assign t[29] = ~(t[47] ^ t[48]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[49] & t[50]);
  assign t[31] = ~(t[51] & t[52]);
  assign t[32] = ~(t[53] | t[54]);
  assign t[33] = ~(t[55] | t[56]);
  assign t[34] = ~(t[142]);
  assign t[35] = ~(t[143]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[59] | t[60]);
  assign t[38] = ~(t[144] | t[61]);
  assign t[39] = t[62] ? x[31] : x[30];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[63] & t[64]);
  assign t[41] = ~(t[65] | t[66]);
  assign t[42] = ~(t[145] | t[67]);
  assign t[43] = ~(t[68] | t[69]);
  assign t[44] = ~(t[70] ^ t[71]);
  assign t[45] = ~(t[72] | t[73]);
  assign t[46] = ~(t[146] | t[74]);
  assign t[47] = ~(t[75] | t[76]);
  assign t[48] = ~(t[77] ^ t[78]);
  assign t[49] = ~(t[79] | t[137]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[80] & t[81]);
  assign t[51] = ~(t[138] | t[82]);
  assign t[52] = t[83] & t[137];
  assign t[53] = ~(t[83] | t[84]);
  assign t[54] = ~(t[83] | t[85]);
  assign t[55] = ~(t[83] | t[86]);
  assign t[56] = ~(t[83] | t[87]);
  assign t[57] = ~(t[147]);
  assign t[58] = ~(t[142] | t[143]);
  assign t[59] = ~(t[148]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[149]);
  assign t[61] = ~(t[88] | t[89]);
  assign t[62] = ~(t[90]);
  assign t[63] = ~(t[20] | t[91]);
  assign t[64] = ~(t[53]);
  assign t[65] = ~(t[150]);
  assign t[66] = ~(t[151]);
  assign t[67] = ~(t[92] | t[93]);
  assign t[68] = ~(t[94] | t[95]);
  assign t[69] = ~(t[152] | t[96]);
  assign t[6] = ~(t[137] & t[138]);
  assign t[70] = t[139] ? x[52] : x[51];
  assign t[71] = ~(t[97] & t[98]);
  assign t[72] = ~(t[153]);
  assign t[73] = ~(t[154]);
  assign t[74] = ~(t[99] | t[100]);
  assign t[75] = ~(t[101] | t[102]);
  assign t[76] = ~(t[155] | t[103]);
  assign t[77] = t[139] ? x[61] : x[60];
  assign t[78] = ~(t[97] & t[104]);
  assign t[79] = ~(t[139]);
  assign t[7] = ~(t[139] & t[140]);
  assign t[80] = ~(t[140] & t[105]);
  assign t[81] = ~(x[4] & t[51]);
  assign t[82] = ~(t[140]);
  assign t[83] = ~(t[79]);
  assign t[84] = t[137] ? t[107] : t[106];
  assign t[85] = t[137] ? t[109] : t[108];
  assign t[86] = t[137] ? t[110] : t[80];
  assign t[87] = t[137] ? t[108] : t[109];
  assign t[88] = ~(t[156]);
  assign t[89] = ~(t[148] | t[149]);
  assign t[8] = ~(t[9] ^ t[11]);
  assign t[90] = ~(t[139]);
  assign t[91] = ~(t[111] & t[112]);
  assign t[92] = ~(t[157]);
  assign t[93] = ~(t[150] | t[151]);
  assign t[94] = ~(t[158]);
  assign t[95] = ~(t[159]);
  assign t[96] = ~(t[113] | t[114]);
  assign t[97] = ~(t[53] | t[115]);
  assign t[98] = ~(t[116] | t[117]);
  assign t[99] = ~(t[160]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = t[0] ? t[1] : t[136];
endmodule

module R1ind186(x, y);
 input [121:0] x;
 output y;

 wire [195:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[105] | t[100]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[149]);
  assign t[105] = ~(t[150]);
  assign t[106] = t[151] ^ x[2];
  assign t[107] = t[152] ^ x[8];
  assign t[108] = t[153] ^ x[11];
  assign t[109] = t[154] ^ x[14];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[155] ^ x[17];
  assign t[111] = t[156] ^ x[22];
  assign t[112] = t[157] ^ x[27];
  assign t[113] = t[158] ^ x[31];
  assign t[114] = t[159] ^ x[33];
  assign t[115] = t[160] ^ x[36];
  assign t[116] = t[161] ^ x[39];
  assign t[117] = t[162] ^ x[44];
  assign t[118] = t[163] ^ x[48];
  assign t[119] = t[164] ^ x[50];
  assign t[11] = t[15] ? x[19] : x[18];
  assign t[120] = t[165] ^ x[53];
  assign t[121] = t[166] ^ x[56];
  assign t[122] = t[167] ^ x[61];
  assign t[123] = t[168] ^ x[65];
  assign t[124] = t[169] ^ x[67];
  assign t[125] = t[170] ^ x[69];
  assign t[126] = t[171] ^ x[71];
  assign t[127] = t[172] ^ x[73];
  assign t[128] = t[173] ^ x[75];
  assign t[129] = t[174] ^ x[77];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[175] ^ x[80];
  assign t[131] = t[176] ^ x[82];
  assign t[132] = t[177] ^ x[84];
  assign t[133] = t[178] ^ x[86];
  assign t[134] = t[179] ^ x[88];
  assign t[135] = t[180] ^ x[90];
  assign t[136] = t[181] ^ x[93];
  assign t[137] = t[182] ^ x[95];
  assign t[138] = t[183] ^ x[97];
  assign t[139] = t[184] ^ x[99];
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = t[185] ^ x[101];
  assign t[141] = t[186] ^ x[103];
  assign t[142] = t[187] ^ x[105];
  assign t[143] = t[188] ^ x[107];
  assign t[144] = t[189] ^ x[109];
  assign t[145] = t[190] ^ x[111];
  assign t[146] = t[191] ^ x[113];
  assign t[147] = t[192] ^ x[115];
  assign t[148] = t[193] ^ x[117];
  assign t[149] = t[194] ^ x[119];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[195] ^ x[121];
  assign t[151] = (x[0] & x[1]);
  assign t[152] = (x[6] & x[7]);
  assign t[153] = (x[9] & x[10]);
  assign t[154] = (x[12] & x[13]);
  assign t[155] = (x[15] & x[16]);
  assign t[156] = (x[20] & x[21]);
  assign t[157] = (x[25] & x[26]);
  assign t[158] = (x[20] & x[30]);
  assign t[159] = (x[20] & x[32]);
  assign t[15] = ~(t[22]);
  assign t[160] = (x[34] & x[35]);
  assign t[161] = (x[37] & x[38]);
  assign t[162] = (x[42] & x[43]);
  assign t[163] = (x[25] & x[47]);
  assign t[164] = (x[25] & x[49]);
  assign t[165] = (x[51] & x[52]);
  assign t[166] = (x[54] & x[55]);
  assign t[167] = (x[59] & x[60]);
  assign t[168] = (x[20] & x[64]);
  assign t[169] = (x[34] & x[66]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[170] = (x[34] & x[68]);
  assign t[171] = (x[37] & x[70]);
  assign t[172] = (x[37] & x[72]);
  assign t[173] = (x[42] & x[74]);
  assign t[174] = (x[42] & x[76]);
  assign t[175] = (x[78] & x[79]);
  assign t[176] = (x[25] & x[81]);
  assign t[177] = (x[51] & x[83]);
  assign t[178] = (x[51] & x[85]);
  assign t[179] = (x[54] & x[87]);
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[180] = (x[54] & x[89]);
  assign t[181] = (x[91] & x[92]);
  assign t[182] = (x[59] & x[94]);
  assign t[183] = (x[59] & x[96]);
  assign t[184] = (x[34] & x[98]);
  assign t[185] = (x[37] & x[100]);
  assign t[186] = (x[42] & x[102]);
  assign t[187] = (x[78] & x[104]);
  assign t[188] = (x[78] & x[106]);
  assign t[189] = (x[51] & x[108]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[190] = (x[54] & x[110]);
  assign t[191] = (x[91] & x[112]);
  assign t[192] = (x[91] & x[114]);
  assign t[193] = (x[59] & x[116]);
  assign t[194] = (x[78] & x[118]);
  assign t[195] = (x[91] & x[120]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[109]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[43] & t[44]);
  assign t[28] = t[45] | t[111];
  assign t[29] = t[15] ? x[24] : x[23];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[39];
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = t[57] | t[112];
  assign t[37] = t[109] ? x[29] : x[28];
  assign t[38] = ~(t[58] & t[59]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[113]);
  assign t[44] = ~(t[114]);
  assign t[45] = ~(t[67] | t[43]);
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = t[70] | t[115];
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = t[73] | t[116];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[74] ? x[41] : x[40];
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = t[77] | t[117];
  assign t[53] = t[74] ? x[46] : x[45];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[118]);
  assign t[56] = ~(t[119]);
  assign t[57] = ~(t[80] | t[55]);
  assign t[58] = ~(t[81] & t[82]);
  assign t[59] = t[83] | t[120];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = t[86] | t[121];
  assign t[62] = t[109] ? x[58] : x[57];
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = t[91] | t[122];
  assign t[66] = t[109] ? x[63] : x[62];
  assign t[67] = ~(t[123]);
  assign t[68] = ~(t[124]);
  assign t[69] = ~(t[125]);
  assign t[6] = ~(t[107] & t[108]);
  assign t[70] = ~(t[92] | t[68]);
  assign t[71] = ~(t[126]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[93] | t[71]);
  assign t[74] = ~(t[22]);
  assign t[75] = ~(t[128]);
  assign t[76] = ~(t[129]);
  assign t[77] = ~(t[94] | t[75]);
  assign t[78] = ~(t[95] & t[96]);
  assign t[79] = t[97] | t[130];
  assign t[7] = ~(t[109] & t[110]);
  assign t[80] = ~(t[131]);
  assign t[81] = ~(t[132]);
  assign t[82] = ~(t[133]);
  assign t[83] = ~(t[98] | t[81]);
  assign t[84] = ~(t[134]);
  assign t[85] = ~(t[135]);
  assign t[86] = ~(t[99] | t[84]);
  assign t[87] = ~(t[100] & t[101]);
  assign t[88] = t[102] | t[136];
  assign t[89] = ~(t[137]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[138]);
  assign t[91] = ~(t[103] | t[89]);
  assign t[92] = ~(t[139]);
  assign t[93] = ~(t[140]);
  assign t[94] = ~(t[141]);
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[104] | t[95]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[145]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[106];
endmodule

module R1ind187(x, y);
 input [121:0] x;
 output y;

 wire [205:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = ~(t[152]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[112] & t[113]);
  assign t[103] = ~(t[143] & t[142]);
  assign t[104] = ~(t[154]);
  assign t[105] = ~(t[145] & t[144]);
  assign t[106] = ~(t[155]);
  assign t[107] = ~(t[156]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[114] & t[115]);
  assign t[10] = x[18] ^ x[19];
  assign t[110] = ~(t[148] & t[147]);
  assign t[111] = ~(t[158]);
  assign t[112] = ~(t[153] & t[152]);
  assign t[113] = ~(t[159]);
  assign t[114] = ~(t[157] & t[156]);
  assign t[115] = ~(t[160]);
  assign t[116] = t[161] ^ x[2];
  assign t[117] = t[162] ^ x[8];
  assign t[118] = t[163] ^ x[11];
  assign t[119] = t[164] ^ x[14];
  assign t[11] = t[15] ? x[18] : x[19];
  assign t[120] = t[165] ^ x[17];
  assign t[121] = t[166] ^ x[22];
  assign t[122] = t[167] ^ x[27];
  assign t[123] = t[168] ^ x[31];
  assign t[124] = t[169] ^ x[33];
  assign t[125] = t[170] ^ x[36];
  assign t[126] = t[171] ^ x[39];
  assign t[127] = t[172] ^ x[44];
  assign t[128] = t[173] ^ x[48];
  assign t[129] = t[174] ^ x[50];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[175] ^ x[53];
  assign t[131] = t[176] ^ x[56];
  assign t[132] = t[177] ^ x[61];
  assign t[133] = t[178] ^ x[65];
  assign t[134] = t[179] ^ x[67];
  assign t[135] = t[180] ^ x[69];
  assign t[136] = t[181] ^ x[71];
  assign t[137] = t[182] ^ x[73];
  assign t[138] = t[183] ^ x[75];
  assign t[139] = t[184] ^ x[77];
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = t[185] ^ x[80];
  assign t[141] = t[186] ^ x[82];
  assign t[142] = t[187] ^ x[84];
  assign t[143] = t[188] ^ x[86];
  assign t[144] = t[189] ^ x[88];
  assign t[145] = t[190] ^ x[90];
  assign t[146] = t[191] ^ x[93];
  assign t[147] = t[192] ^ x[95];
  assign t[148] = t[193] ^ x[97];
  assign t[149] = t[194] ^ x[99];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[195] ^ x[101];
  assign t[151] = t[196] ^ x[103];
  assign t[152] = t[197] ^ x[105];
  assign t[153] = t[198] ^ x[107];
  assign t[154] = t[199] ^ x[109];
  assign t[155] = t[200] ^ x[111];
  assign t[156] = t[201] ^ x[113];
  assign t[157] = t[202] ^ x[115];
  assign t[158] = t[203] ^ x[117];
  assign t[159] = t[204] ^ x[119];
  assign t[15] = ~(t[22]);
  assign t[160] = t[205] ^ x[121];
  assign t[161] = (x[0] & x[1]);
  assign t[162] = (x[6] & x[7]);
  assign t[163] = (x[9] & x[10]);
  assign t[164] = (x[12] & x[13]);
  assign t[165] = (x[15] & x[16]);
  assign t[166] = (x[20] & x[21]);
  assign t[167] = (x[25] & x[26]);
  assign t[168] = (x[20] & x[30]);
  assign t[169] = (x[20] & x[32]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[170] = (x[34] & x[35]);
  assign t[171] = (x[37] & x[38]);
  assign t[172] = (x[42] & x[43]);
  assign t[173] = (x[25] & x[47]);
  assign t[174] = (x[25] & x[49]);
  assign t[175] = (x[51] & x[52]);
  assign t[176] = (x[54] & x[55]);
  assign t[177] = (x[59] & x[60]);
  assign t[178] = (x[20] & x[64]);
  assign t[179] = (x[34] & x[66]);
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[180] = (x[34] & x[68]);
  assign t[181] = (x[37] & x[70]);
  assign t[182] = (x[37] & x[72]);
  assign t[183] = (x[42] & x[74]);
  assign t[184] = (x[42] & x[76]);
  assign t[185] = (x[78] & x[79]);
  assign t[186] = (x[25] & x[81]);
  assign t[187] = (x[51] & x[83]);
  assign t[188] = (x[51] & x[85]);
  assign t[189] = (x[54] & x[87]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[190] = (x[54] & x[89]);
  assign t[191] = (x[91] & x[92]);
  assign t[192] = (x[59] & x[94]);
  assign t[193] = (x[59] & x[96]);
  assign t[194] = (x[34] & x[98]);
  assign t[195] = (x[37] & x[100]);
  assign t[196] = (x[42] & x[102]);
  assign t[197] = (x[78] & x[104]);
  assign t[198] = (x[78] & x[106]);
  assign t[199] = (x[51] & x[108]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[200] = (x[54] & x[110]);
  assign t[201] = (x[91] & x[112]);
  assign t[202] = (x[91] & x[114]);
  assign t[203] = (x[59] & x[116]);
  assign t[204] = (x[78] & x[118]);
  assign t[205] = (x[91] & x[120]);
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[119]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[43] & t[44]);
  assign t[28] = ~(t[45] & t[121]);
  assign t[29] = t[46] ? x[24] : x[23];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = ~(t[49] & t[50]);
  assign t[32] = t[51] ^ t[39];
  assign t[33] = ~(t[52] & t[53]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = ~(t[56] & t[57]);
  assign t[36] = ~(t[58] & t[122]);
  assign t[37] = t[119] ? x[29] : x[28];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = ~(t[61] & t[62]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[63] ^ t[64];
  assign t[41] = ~(t[65] & t[66]);
  assign t[42] = t[67] ^ t[41];
  assign t[43] = ~(t[123]);
  assign t[44] = ~(t[124]);
  assign t[45] = ~(t[68] & t[69]);
  assign t[46] = ~(t[22]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[125]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[75] & t[126]);
  assign t[51] = t[15] ? x[41] : x[40];
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = ~(t[78] & t[127]);
  assign t[54] = t[15] ? x[46] : x[45];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[128]);
  assign t[57] = ~(t[129]);
  assign t[58] = ~(t[81] & t[82]);
  assign t[59] = ~(t[83] & t[84]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[85] & t[130]);
  assign t[61] = ~(t[86] & t[87]);
  assign t[62] = ~(t[88] & t[131]);
  assign t[63] = t[119] ? x[58] : x[57];
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[92]);
  assign t[66] = ~(t[93] & t[132]);
  assign t[67] = t[119] ? x[63] : x[62];
  assign t[68] = ~(t[124] & t[123]);
  assign t[69] = ~(t[133]);
  assign t[6] = ~(t[117] & t[118]);
  assign t[70] = ~(t[134]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[94] & t[95]);
  assign t[73] = ~(t[136]);
  assign t[74] = ~(t[137]);
  assign t[75] = ~(t[96] & t[97]);
  assign t[76] = ~(t[138]);
  assign t[77] = ~(t[139]);
  assign t[78] = ~(t[98] & t[99]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = ~(t[119] & t[120]);
  assign t[80] = ~(t[102] & t[140]);
  assign t[81] = ~(t[129] & t[128]);
  assign t[82] = ~(t[141]);
  assign t[83] = ~(t[142]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[103] & t[104]);
  assign t[86] = ~(t[144]);
  assign t[87] = ~(t[145]);
  assign t[88] = ~(t[105] & t[106]);
  assign t[89] = ~(t[107] & t[108]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[109] & t[146]);
  assign t[91] = ~(t[147]);
  assign t[92] = ~(t[148]);
  assign t[93] = ~(t[110] & t[111]);
  assign t[94] = ~(t[135] & t[134]);
  assign t[95] = ~(t[149]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[150]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[151]);
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[116];
endmodule

module R1ind188(x, y);
 input [101:0] x;
 output y;

 wire [166:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[135] ^ x[14];
  assign t[101] = t[136] ^ x[17];
  assign t[102] = t[137] ^ x[22];
  assign t[103] = t[138] ^ x[24];
  assign t[104] = t[139] ^ x[29];
  assign t[105] = t[140] ^ x[31];
  assign t[106] = t[141] ^ x[35];
  assign t[107] = t[142] ^ x[38];
  assign t[108] = t[143] ^ x[40];
  assign t[109] = t[144] ^ x[43];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[145] ^ x[45];
  assign t[111] = t[146] ^ x[50];
  assign t[112] = t[147] ^ x[52];
  assign t[113] = t[148] ^ x[56];
  assign t[114] = t[149] ^ x[59];
  assign t[115] = t[150] ^ x[61];
  assign t[116] = t[151] ^ x[64];
  assign t[117] = t[152] ^ x[66];
  assign t[118] = t[153] ^ x[71];
  assign t[119] = t[154] ^ x[73];
  assign t[11] = t[15] ? x[18] : x[19];
  assign t[120] = t[155] ^ x[77];
  assign t[121] = t[156] ^ x[79];
  assign t[122] = t[157] ^ x[81];
  assign t[123] = t[158] ^ x[84];
  assign t[124] = t[159] ^ x[86];
  assign t[125] = t[160] ^ x[88];
  assign t[126] = t[161] ^ x[90];
  assign t[127] = t[162] ^ x[92];
  assign t[128] = t[163] ^ x[95];
  assign t[129] = t[164] ^ x[97];
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = t[165] ^ x[99];
  assign t[131] = t[166] ^ x[101];
  assign t[132] = (x[0] & x[1]);
  assign t[133] = (x[6] & x[7]);
  assign t[134] = (x[9] & x[10]);
  assign t[135] = (x[12] & x[13]);
  assign t[136] = (x[15] & x[16]);
  assign t[137] = (x[20] & x[21]);
  assign t[138] = (x[20] & x[23]);
  assign t[139] = (x[27] & x[28]);
  assign t[13] = x[4] ? t[19] : t[18];
  assign t[140] = (x[27] & x[30]);
  assign t[141] = (x[20] & x[34]);
  assign t[142] = (x[36] & x[37]);
  assign t[143] = (x[36] & x[39]);
  assign t[144] = (x[41] & x[42]);
  assign t[145] = (x[41] & x[44]);
  assign t[146] = (x[48] & x[49]);
  assign t[147] = (x[48] & x[51]);
  assign t[148] = (x[27] & x[55]);
  assign t[149] = (x[57] & x[58]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (x[57] & x[60]);
  assign t[151] = (x[62] & x[63]);
  assign t[152] = (x[62] & x[65]);
  assign t[153] = (x[69] & x[70]);
  assign t[154] = (x[69] & x[72]);
  assign t[155] = (x[36] & x[76]);
  assign t[156] = (x[41] & x[78]);
  assign t[157] = (x[48] & x[80]);
  assign t[158] = (x[82] & x[83]);
  assign t[159] = (x[82] & x[85]);
  assign t[15] = ~(t[22]);
  assign t[160] = (x[57] & x[87]);
  assign t[161] = (x[62] & x[89]);
  assign t[162] = (x[69] & x[91]);
  assign t[163] = (x[93] & x[94]);
  assign t[164] = (x[93] & x[96]);
  assign t[165] = (x[82] & x[98]);
  assign t[166] = (x[93] & x[100]);
  assign t[16] = x[4] ? t[24] : t[23];
  assign t[17] = ~(t[25] ^ t[26]);
  assign t[18] = ~(t[27] & t[28]);
  assign t[19] = t[29] ^ t[30];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[32] : t[31];
  assign t[21] = x[4] ? t[34] : t[33];
  assign t[22] = ~(t[100]);
  assign t[23] = ~(t[35] & t[36]);
  assign t[24] = t[37] ^ t[38];
  assign t[25] = x[4] ? t[40] : t[39];
  assign t[26] = x[4] ? t[42] : t[41];
  assign t[27] = ~(t[102] & t[43]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[29] = t[45] ? x[26] : x[25];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[41];
  assign t[33] = ~(t[51] & t[52]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = ~(t[104] & t[55]);
  assign t[36] = ~(t[105] & t[56]);
  assign t[37] = t[100] ? x[33] : x[32];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = ~(x[3]);
  assign t[40] = t[61] ^ t[39];
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[106]);
  assign t[44] = ~(t[106] & t[66]);
  assign t[45] = ~(t[22]);
  assign t[46] = ~(t[107] & t[67]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[71] ? x[47] : x[46];
  assign t[51] = ~(t[111] & t[72]);
  assign t[52] = ~(t[112] & t[73]);
  assign t[53] = t[71] ? x[54] : x[53];
  assign t[54] = ~(t[74] & t[75]);
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[113] & t[76]);
  assign t[57] = ~(t[114] & t[77]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = t[100] ? x[68] : x[67];
  assign t[62] = ~(t[118] & t[81]);
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = t[100] ? x[75] : x[74];
  assign t[65] = ~(t[83] & t[84]);
  assign t[66] = ~(t[102]);
  assign t[67] = ~(t[120]);
  assign t[68] = ~(t[120] & t[85]);
  assign t[69] = ~(t[121]);
  assign t[6] = ~(t[98] & t[99]);
  assign t[70] = ~(t[121] & t[86]);
  assign t[71] = ~(t[22]);
  assign t[72] = ~(t[122]);
  assign t[73] = ~(t[122] & t[87]);
  assign t[74] = ~(t[123] & t[88]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[104]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[125] & t[90]);
  assign t[79] = ~(t[126]);
  assign t[7] = ~(t[100] & t[101]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[127] & t[92]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[107]);
  assign t[86] = ~(t[109]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[130]);
  assign t[89] = ~(t[130] & t[95]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[114]);
  assign t[91] = ~(t[116]);
  assign t[92] = ~(t[118]);
  assign t[93] = ~(t[131]);
  assign t[94] = ~(t[131] & t[96]);
  assign t[95] = ~(t[123]);
  assign t[96] = ~(t[128]);
  assign t[97] = t[132] ^ x[2];
  assign t[98] = t[133] ^ x[8];
  assign t[99] = t[134] ^ x[11];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[97];
endmodule

module R1ind189(x, y);
 input [121:0] x;
 output y;

 wire [293:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[145] ? x[70] : x[69];
  assign t[101] = ~(t[146] & t[82]);
  assign t[102] = ~(t[227]);
  assign t[103] = ~(t[228]);
  assign t[104] = ~(t[147] | t[148]);
  assign t[105] = t[145] ? x[76] : x[75];
  assign t[106] = ~(t[149] & t[150]);
  assign t[107] = ~(t[229]);
  assign t[108] = ~(t[216] | t[217]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(x[3]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[151] | t[152]);
  assign t[112] = ~(t[153] | t[154]);
  assign t[113] = ~(t[232]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[155] | t[156]);
  assign t[116] = ~(t[157] | t[158]);
  assign t[117] = ~(t[234] | t[159]);
  assign t[118] = t[92] ? x[91] : x[90];
  assign t[119] = ~(t[160] & t[161]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[235]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[162] | t[163]);
  assign t[123] = t[207] ? x[97] : x[96];
  assign t[124] = t[164] | t[165];
  assign t[125] = ~(t[166] & t[208]);
  assign t[126] = ~(t[167] & t[168]);
  assign t[127] = ~(t[79] | t[169]);
  assign t[128] = ~(t[79] | t[170]);
  assign t[129] = t[208] & t[171];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = t[167] | t[166];
  assign t[131] = ~(x[4] & t[172]);
  assign t[132] = ~(t[173] & t[168]);
  assign t[133] = t[205] ? t[175] : t[174];
  assign t[134] = ~(t[171] & t[176]);
  assign t[135] = ~(t[237]);
  assign t[136] = ~(t[222] | t[223]);
  assign t[137] = ~(t[207]);
  assign t[138] = ~(t[112]);
  assign t[139] = ~(t[79] | t[177]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[238]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[239]);
  assign t[143] = ~(t[240]);
  assign t[144] = ~(t[178] | t[179]);
  assign t[145] = ~(t[137]);
  assign t[146] = ~(t[164] | t[180]);
  assign t[147] = ~(t[241]);
  assign t[148] = ~(t[227] | t[228]);
  assign t[149] = ~(t[127] | t[181]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[182] & t[183]);
  assign t[151] = ~(t[242]);
  assign t[152] = ~(t[230] | t[231]);
  assign t[153] = ~(t[79] | t[184]);
  assign t[154] = ~(t[79] | t[185]);
  assign t[155] = ~(t[243]);
  assign t[156] = ~(t[232] | t[233]);
  assign t[157] = ~(t[244]);
  assign t[158] = ~(t[245]);
  assign t[159] = ~(t[186] | t[187]);
  assign t[15] = ~(t[205] & t[206]);
  assign t[160] = ~(t[164] | t[188]);
  assign t[161] = ~(t[47]);
  assign t[162] = ~(t[246]);
  assign t[163] = ~(t[235] | t[236]);
  assign t[164] = ~(t[134] & t[150]);
  assign t[165] = ~(t[189] & t[190]);
  assign t[166] = x[4] & t[206];
  assign t[167] = ~(x[4] | t[206]);
  assign t[168] = ~(t[208]);
  assign t[169] = t[205] ? t[125] : t[126];
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = t[205] ? t[131] : t[191];
  assign t[171] = ~(t[83] | t[205]);
  assign t[172] = ~(t[206] | t[208]);
  assign t[173] = ~(x[4] | t[192]);
  assign t[174] = ~(t[166] & t[168]);
  assign t[175] = ~(t[167] & t[208]);
  assign t[176] = ~(t[191] & t[193]);
  assign t[177] = t[205] ? t[191] : t[131];
  assign t[178] = ~(t[247]);
  assign t[179] = ~(t[239] | t[240]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = t[139] | t[85];
  assign t[181] = ~(t[194] & t[195]);
  assign t[182] = ~(t[206] | t[168]);
  assign t[183] = t[79] & t[205];
  assign t[184] = t[205] ? t[193] : t[132];
  assign t[185] = t[205] ? t[174] : t[175];
  assign t[186] = ~(t[248]);
  assign t[187] = ~(t[244] | t[245]);
  assign t[188] = ~(t[196] & t[197]);
  assign t[189] = ~(t[47] | t[85]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = ~(t[128] | t[154]);
  assign t[191] = ~(t[208] & t[173]);
  assign t[192] = ~(t[206]);
  assign t[193] = ~(x[4] & t[182]);
  assign t[194] = ~(t[198] | t[199]);
  assign t[195] = ~(t[83] & t[200]);
  assign t[196] = ~(t[49]);
  assign t[197] = t[83] | t[201];
  assign t[198] = ~(t[83] | t[202]);
  assign t[199] = ~(t[79] | t[203]);
  assign t[19] = t[207] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = ~(t[131] & t[191]);
  assign t[201] = t[205] ? t[131] : t[132];
  assign t[202] = t[205] ? t[126] : t[174];
  assign t[203] = t[205] ? t[132] : t[193];
  assign t[204] = t[249] ^ x[2];
  assign t[205] = t[250] ^ x[10];
  assign t[206] = t[251] ^ x[13];
  assign t[207] = t[252] ^ x[16];
  assign t[208] = t[253] ^ x[19];
  assign t[209] = t[254] ^ x[22];
  assign t[20] = ~(t[29] & t[30]);
  assign t[210] = t[255] ^ x[25];
  assign t[211] = t[256] ^ x[27];
  assign t[212] = t[257] ^ x[29];
  assign t[213] = t[258] ^ x[32];
  assign t[214] = t[259] ^ x[37];
  assign t[215] = t[260] ^ x[40];
  assign t[216] = t[261] ^ x[42];
  assign t[217] = t[262] ^ x[44];
  assign t[218] = t[263] ^ x[47];
  assign t[219] = t[264] ^ x[52];
  assign t[21] = ~(t[31] | t[32]);
  assign t[220] = t[265] ^ x[55];
  assign t[221] = t[266] ^ x[57];
  assign t[222] = t[267] ^ x[59];
  assign t[223] = t[268] ^ x[61];
  assign t[224] = t[269] ^ x[63];
  assign t[225] = t[270] ^ x[65];
  assign t[226] = t[271] ^ x[68];
  assign t[227] = t[272] ^ x[72];
  assign t[228] = t[273] ^ x[74];
  assign t[229] = t[274] ^ x[78];
  assign t[22] = ~(t[33] ^ t[34]);
  assign t[230] = t[275] ^ x[80];
  assign t[231] = t[276] ^ x[82];
  assign t[232] = t[277] ^ x[84];
  assign t[233] = t[278] ^ x[86];
  assign t[234] = t[279] ^ x[89];
  assign t[235] = t[280] ^ x[93];
  assign t[236] = t[281] ^ x[95];
  assign t[237] = t[282] ^ x[99];
  assign t[238] = t[283] ^ x[101];
  assign t[239] = t[284] ^ x[103];
  assign t[23] = x[4] ? t[36] : t[35];
  assign t[240] = t[285] ^ x[105];
  assign t[241] = t[286] ^ x[107];
  assign t[242] = t[287] ^ x[109];
  assign t[243] = t[288] ^ x[111];
  assign t[244] = t[289] ^ x[113];
  assign t[245] = t[290] ^ x[115];
  assign t[246] = t[291] ^ x[117];
  assign t[247] = t[292] ^ x[119];
  assign t[248] = t[293] ^ x[121];
  assign t[249] = (x[0] & x[1]);
  assign t[24] = x[4] ? t[38] : t[37];
  assign t[250] = (x[8] & x[9]);
  assign t[251] = (x[11] & x[12]);
  assign t[252] = (x[14] & x[15]);
  assign t[253] = (x[17] & x[18]);
  assign t[254] = (x[20] & x[21]);
  assign t[255] = (x[23] & x[24]);
  assign t[256] = (x[20] & x[26]);
  assign t[257] = (x[20] & x[28]);
  assign t[258] = (x[30] & x[31]);
  assign t[259] = (x[35] & x[36]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[260] = (x[38] & x[39]);
  assign t[261] = (x[23] & x[41]);
  assign t[262] = (x[23] & x[43]);
  assign t[263] = (x[45] & x[46]);
  assign t[264] = (x[50] & x[51]);
  assign t[265] = (x[53] & x[54]);
  assign t[266] = (x[20] & x[56]);
  assign t[267] = (x[30] & x[58]);
  assign t[268] = (x[30] & x[60]);
  assign t[269] = (x[35] & x[62]);
  assign t[26] = ~(t[41] ^ t[42]);
  assign t[270] = (x[35] & x[64]);
  assign t[271] = (x[66] & x[67]);
  assign t[272] = (x[38] & x[71]);
  assign t[273] = (x[38] & x[73]);
  assign t[274] = (x[23] & x[77]);
  assign t[275] = (x[45] & x[79]);
  assign t[276] = (x[45] & x[81]);
  assign t[277] = (x[50] & x[83]);
  assign t[278] = (x[50] & x[85]);
  assign t[279] = (x[87] & x[88]);
  assign t[27] = x[4] ? t[44] : t[43];
  assign t[280] = (x[53] & x[92]);
  assign t[281] = (x[53] & x[94]);
  assign t[282] = (x[30] & x[98]);
  assign t[283] = (x[35] & x[100]);
  assign t[284] = (x[66] & x[102]);
  assign t[285] = (x[66] & x[104]);
  assign t[286] = (x[38] & x[106]);
  assign t[287] = (x[45] & x[108]);
  assign t[288] = (x[50] & x[110]);
  assign t[289] = (x[87] & x[112]);
  assign t[28] = x[4] ? t[46] : t[45];
  assign t[290] = (x[87] & x[114]);
  assign t[291] = (x[53] & x[116]);
  assign t[292] = (x[66] & x[118]);
  assign t[293] = (x[87] & x[120]);
  assign t[29] = ~(t[47] | t[48]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[49] | t[50]);
  assign t[31] = ~(t[51] | t[52]);
  assign t[32] = ~(t[209] | t[53]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[34] = ~(t[56] ^ t[57]);
  assign t[35] = ~(t[58] | t[59]);
  assign t[36] = ~(t[60] ^ t[61]);
  assign t[37] = ~(t[62] | t[63]);
  assign t[38] = ~(t[43] ^ t[64]);
  assign t[39] = ~(t[65] | t[66]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[210] | t[67]);
  assign t[41] = ~(t[68] | t[69]);
  assign t[42] = ~(t[70] ^ t[71]);
  assign t[43] = ~(t[72] | t[73]);
  assign t[44] = ~(t[74] ^ t[75]);
  assign t[45] = ~(t[76] | t[77]);
  assign t[46] = ~(t[45] ^ t[78]);
  assign t[47] = ~(t[79] | t[80]);
  assign t[48] = ~(t[81] & t[82]);
  assign t[49] = ~(t[83] | t[84]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[85] | t[86];
  assign t[51] = ~(t[211]);
  assign t[52] = ~(t[212]);
  assign t[53] = ~(t[87] | t[88]);
  assign t[54] = ~(t[89] | t[90]);
  assign t[55] = ~(t[213] | t[91]);
  assign t[56] = t[92] ? x[34] : x[33];
  assign t[57] = ~(t[93] & t[94]);
  assign t[58] = ~(t[95] | t[96]);
  assign t[59] = ~(t[214] | t[97]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[98] | t[99]);
  assign t[61] = ~(t[100] ^ t[101]);
  assign t[62] = ~(t[102] | t[103]);
  assign t[63] = ~(t[215] | t[104]);
  assign t[64] = ~(t[105] ^ t[106]);
  assign t[65] = ~(t[216]);
  assign t[66] = ~(t[217]);
  assign t[67] = ~(t[107] | t[108]);
  assign t[68] = ~(t[109] | t[110]);
  assign t[69] = ~(t[218] | t[111]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[207] ? x[49] : x[48];
  assign t[71] = ~(t[29] & t[112]);
  assign t[72] = ~(t[113] | t[114]);
  assign t[73] = ~(t[219] | t[115]);
  assign t[74] = ~(t[116] | t[117]);
  assign t[75] = ~(t[118] ^ t[119]);
  assign t[76] = ~(t[120] | t[121]);
  assign t[77] = ~(t[220] | t[122]);
  assign t[78] = ~(t[123] ^ t[124]);
  assign t[79] = ~(t[83]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[205] ? t[126] : t[125];
  assign t[81] = ~(t[127] | t[128]);
  assign t[82] = ~(t[129] & t[130]);
  assign t[83] = ~(t[207]);
  assign t[84] = t[205] ? t[132] : t[131];
  assign t[85] = ~(t[79] | t[133]);
  assign t[86] = ~(t[134]);
  assign t[87] = ~(t[221]);
  assign t[88] = ~(t[211] | t[212]);
  assign t[89] = ~(t[222]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[223]);
  assign t[91] = ~(t[135] | t[136]);
  assign t[92] = ~(t[137]);
  assign t[93] = ~(t[127]);
  assign t[94] = ~(t[138] | t[139]);
  assign t[95] = ~(t[224]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[140] | t[141]);
  assign t[98] = ~(t[142] | t[143]);
  assign t[99] = ~(t[226] | t[144]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[204];
endmodule

module R1ind190(x, y);
 input [112:0] x;
 output y;

 wire [180:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[141] ^ x[8];
  assign t[101] = t[142] ^ x[11];
  assign t[102] = t[143] ^ x[14];
  assign t[103] = t[144] ^ x[17];
  assign t[104] = t[145] ^ x[22];
  assign t[105] = t[146] ^ x[27];
  assign t[106] = t[147] ^ x[31];
  assign t[107] = t[148] ^ x[33];
  assign t[108] = t[149] ^ x[36];
  assign t[109] = t[150] ^ x[41];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[151] ^ x[45];
  assign t[111] = t[152] ^ x[47];
  assign t[112] = t[153] ^ x[50];
  assign t[113] = t[154] ^ x[53];
  assign t[114] = t[155] ^ x[58];
  assign t[115] = t[156] ^ x[62];
  assign t[116] = t[157] ^ x[64];
  assign t[117] = t[158] ^ x[66];
  assign t[118] = t[159] ^ x[68];
  assign t[119] = t[160] ^ x[70];
  assign t[11] = t[102] ? x[18] : x[19];
  assign t[120] = t[161] ^ x[73];
  assign t[121] = t[162] ^ x[75];
  assign t[122] = t[163] ^ x[77];
  assign t[123] = t[164] ^ x[79];
  assign t[124] = t[165] ^ x[81];
  assign t[125] = t[166] ^ x[83];
  assign t[126] = t[167] ^ x[86];
  assign t[127] = t[168] ^ x[88];
  assign t[128] = t[169] ^ x[90];
  assign t[129] = t[170] ^ x[92];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = t[171] ^ x[94];
  assign t[131] = t[172] ^ x[96];
  assign t[132] = t[173] ^ x[98];
  assign t[133] = t[174] ^ x[100];
  assign t[134] = t[175] ^ x[102];
  assign t[135] = t[176] ^ x[104];
  assign t[136] = t[177] ^ x[106];
  assign t[137] = t[178] ^ x[108];
  assign t[138] = t[179] ^ x[110];
  assign t[139] = t[180] ^ x[112];
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (x[0] & x[1]);
  assign t[141] = (x[6] & x[7]);
  assign t[142] = (x[9] & x[10]);
  assign t[143] = (x[12] & x[13]);
  assign t[144] = (x[15] & x[16]);
  assign t[145] = (x[20] & x[21]);
  assign t[146] = (x[25] & x[26]);
  assign t[147] = (x[20] & x[30]);
  assign t[148] = (x[20] & x[32]);
  assign t[149] = (x[34] & x[35]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[39] & x[40]);
  assign t[151] = (x[25] & x[44]);
  assign t[152] = (x[25] & x[46]);
  assign t[153] = (x[48] & x[49]);
  assign t[154] = (x[51] & x[52]);
  assign t[155] = (x[56] & x[57]);
  assign t[156] = (x[20] & x[61]);
  assign t[157] = (x[34] & x[63]);
  assign t[158] = (x[34] & x[65]);
  assign t[159] = (x[39] & x[67]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[160] = (x[39] & x[69]);
  assign t[161] = (x[71] & x[72]);
  assign t[162] = (x[25] & x[74]);
  assign t[163] = (x[48] & x[76]);
  assign t[164] = (x[48] & x[78]);
  assign t[165] = (x[51] & x[80]);
  assign t[166] = (x[51] & x[82]);
  assign t[167] = (x[84] & x[85]);
  assign t[168] = (x[56] & x[87]);
  assign t[169] = (x[56] & x[89]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (x[34] & x[91]);
  assign t[171] = (x[39] & x[93]);
  assign t[172] = (x[71] & x[95]);
  assign t[173] = (x[71] & x[97]);
  assign t[174] = (x[48] & x[99]);
  assign t[175] = (x[51] & x[101]);
  assign t[176] = (x[84] & x[103]);
  assign t[177] = (x[84] & x[105]);
  assign t[178] = (x[56] & x[107]);
  assign t[179] = (x[71] & x[109]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[180] = (x[84] & x[111]);
  assign t[18] = t[27] ^ t[21];
  assign t[19] = x[4] ? t[29] : t[28];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[21] = ~(t[32] & t[33]);
  assign t[22] = t[34] ^ t[35];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[40] & t[41]);
  assign t[26] = t[42] | t[104];
  assign t[27] = t[43] ? x[24] : x[23];
  assign t[28] = ~(t[44] & t[45]);
  assign t[29] = t[46] ^ t[28];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = t[49] ^ t[50];
  assign t[32] = ~(t[51] & t[52]);
  assign t[33] = t[53] | t[105];
  assign t[34] = t[54] ? x[29] : x[28];
  assign t[35] = ~(t[55] & t[56]);
  assign t[36] = ~(t[57] & t[58]);
  assign t[37] = t[59] ^ t[60];
  assign t[38] = ~(t[61] & t[62]);
  assign t[39] = t[63] ^ t[38];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[106]);
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[64] | t[40]);
  assign t[43] = ~(t[65]);
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] | t[108];
  assign t[46] = t[43] ? x[38] : x[37];
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = t[71] | t[109];
  assign t[49] = t[43] ? x[43] : x[42];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = ~(t[110]);
  assign t[52] = ~(t[111]);
  assign t[53] = ~(t[74] | t[51]);
  assign t[54] = ~(t[65]);
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = t[77] | t[112];
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = t[80] | t[113];
  assign t[59] = t[102] ? x[55] : x[54];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = t[85] | t[114];
  assign t[63] = t[102] ? x[60] : x[59];
  assign t[64] = ~(t[115]);
  assign t[65] = ~(t[102]);
  assign t[66] = ~(t[116]);
  assign t[67] = ~(t[117]);
  assign t[68] = ~(t[86] | t[66]);
  assign t[69] = ~(t[118]);
  assign t[6] = ~(t[100] & t[101]);
  assign t[70] = ~(t[119]);
  assign t[71] = ~(t[87] | t[69]);
  assign t[72] = ~(t[88] & t[89]);
  assign t[73] = t[90] | t[120];
  assign t[74] = ~(t[121]);
  assign t[75] = ~(t[122]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[91] | t[75]);
  assign t[78] = ~(t[124]);
  assign t[79] = ~(t[125]);
  assign t[7] = ~(t[102] & t[103]);
  assign t[80] = ~(t[92] | t[78]);
  assign t[81] = ~(t[93] & t[94]);
  assign t[82] = t[95] | t[126];
  assign t[83] = ~(t[127]);
  assign t[84] = ~(t[128]);
  assign t[85] = ~(t[96] | t[83]);
  assign t[86] = ~(t[129]);
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = ~(t[97] | t[88]);
  assign t[91] = ~(t[133]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[98] | t[93]);
  assign t[96] = ~(t[137]);
  assign t[97] = ~(t[138]);
  assign t[98] = ~(t[139]);
  assign t[99] = t[140] ^ x[2];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[99];
endmodule

module R1ind191(x, y);
 input [112:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[145]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[108] & t[109]);
  assign t[104] = ~(t[139] & t[138]);
  assign t[105] = ~(t[148]);
  assign t[106] = ~(t[143] & t[142]);
  assign t[107] = ~(t[149]);
  assign t[108] = ~(t[147] & t[146]);
  assign t[109] = ~(t[150]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[151] ^ x[2];
  assign t[111] = t[152] ^ x[10];
  assign t[112] = t[153] ^ x[13];
  assign t[113] = t[154] ^ x[16];
  assign t[114] = t[155] ^ x[19];
  assign t[115] = t[156] ^ x[22];
  assign t[116] = t[157] ^ x[27];
  assign t[117] = t[158] ^ x[31];
  assign t[118] = t[159] ^ x[33];
  assign t[119] = t[160] ^ x[36];
  assign t[11] = t[111] ? x[6] : x[7];
  assign t[120] = t[161] ^ x[41];
  assign t[121] = t[162] ^ x[45];
  assign t[122] = t[163] ^ x[47];
  assign t[123] = t[164] ^ x[50];
  assign t[124] = t[165] ^ x[53];
  assign t[125] = t[166] ^ x[58];
  assign t[126] = t[167] ^ x[62];
  assign t[127] = t[168] ^ x[64];
  assign t[128] = t[169] ^ x[66];
  assign t[129] = t[170] ^ x[68];
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[130] = t[171] ^ x[70];
  assign t[131] = t[172] ^ x[73];
  assign t[132] = t[173] ^ x[75];
  assign t[133] = t[174] ^ x[77];
  assign t[134] = t[175] ^ x[79];
  assign t[135] = t[176] ^ x[81];
  assign t[136] = t[177] ^ x[83];
  assign t[137] = t[178] ^ x[86];
  assign t[138] = t[179] ^ x[88];
  assign t[139] = t[180] ^ x[90];
  assign t[13] = x[4] ? t[20] : t[19];
  assign t[140] = t[181] ^ x[92];
  assign t[141] = t[182] ^ x[94];
  assign t[142] = t[183] ^ x[96];
  assign t[143] = t[184] ^ x[98];
  assign t[144] = t[185] ^ x[100];
  assign t[145] = t[186] ^ x[102];
  assign t[146] = t[187] ^ x[104];
  assign t[147] = t[188] ^ x[106];
  assign t[148] = t[189] ^ x[108];
  assign t[149] = t[190] ^ x[110];
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = t[191] ^ x[112];
  assign t[151] = (x[0] & x[1]);
  assign t[152] = (x[8] & x[9]);
  assign t[153] = (x[11] & x[12]);
  assign t[154] = (x[14] & x[15]);
  assign t[155] = (x[17] & x[18]);
  assign t[156] = (x[20] & x[21]);
  assign t[157] = (x[25] & x[26]);
  assign t[158] = (x[20] & x[30]);
  assign t[159] = (x[20] & x[32]);
  assign t[15] = ~(t[112] & t[113]);
  assign t[160] = (x[34] & x[35]);
  assign t[161] = (x[39] & x[40]);
  assign t[162] = (x[25] & x[44]);
  assign t[163] = (x[25] & x[46]);
  assign t[164] = (x[48] & x[49]);
  assign t[165] = (x[51] & x[52]);
  assign t[166] = (x[56] & x[57]);
  assign t[167] = (x[20] & x[61]);
  assign t[168] = (x[34] & x[63]);
  assign t[169] = (x[34] & x[65]);
  assign t[16] = ~(t[111] & t[114]);
  assign t[170] = (x[39] & x[67]);
  assign t[171] = (x[39] & x[69]);
  assign t[172] = (x[71] & x[72]);
  assign t[173] = (x[25] & x[74]);
  assign t[174] = (x[48] & x[76]);
  assign t[175] = (x[48] & x[78]);
  assign t[176] = (x[51] & x[80]);
  assign t[177] = (x[51] & x[82]);
  assign t[178] = (x[84] & x[85]);
  assign t[179] = (x[56] & x[87]);
  assign t[17] = x[4] ? t[24] : t[23];
  assign t[180] = (x[56] & x[89]);
  assign t[181] = (x[34] & x[91]);
  assign t[182] = (x[39] & x[93]);
  assign t[183] = (x[71] & x[95]);
  assign t[184] = (x[71] & x[97]);
  assign t[185] = (x[48] & x[99]);
  assign t[186] = (x[51] & x[101]);
  assign t[187] = (x[84] & x[103]);
  assign t[188] = (x[84] & x[105]);
  assign t[189] = (x[56] & x[107]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[190] = (x[71] & x[109]);
  assign t[191] = (x[84] & x[111]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[29] ^ t[23];
  assign t[21] = x[4] ? t[31] : t[30];
  assign t[22] = x[4] ? t[33] : t[32];
  assign t[23] = ~(t[34] & t[35]);
  assign t[24] = t[36] ^ t[37];
  assign t[25] = x[4] ? t[39] : t[38];
  assign t[26] = x[4] ? t[41] : t[40];
  assign t[27] = ~(t[42] & t[43]);
  assign t[28] = ~(t[44] & t[115]);
  assign t[29] = t[45] ? x[24] : x[23];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = t[48] ^ t[30];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = t[51] ^ t[52];
  assign t[34] = ~(t[53] & t[54]);
  assign t[35] = ~(t[55] & t[116]);
  assign t[36] = t[56] ? x[29] : x[28];
  assign t[37] = ~(t[57] & t[58]);
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[63] & t[64]);
  assign t[41] = t[65] ^ t[40];
  assign t[42] = ~(t[117]);
  assign t[43] = ~(t[118]);
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = ~(t[68]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[71] & t[119]);
  assign t[48] = t[45] ? x[38] : x[37];
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[74] & t[120]);
  assign t[51] = t[45] ? x[43] : x[42];
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = ~(t[121]);
  assign t[54] = ~(t[122]);
  assign t[55] = ~(t[77] & t[78]);
  assign t[56] = ~(t[68]);
  assign t[57] = ~(t[79] & t[80]);
  assign t[58] = ~(t[81] & t[123]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[84] & t[124]);
  assign t[61] = t[111] ? x[55] : x[54];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = ~(t[89] & t[125]);
  assign t[65] = t[111] ? x[60] : x[59];
  assign t[66] = ~(t[118] & t[117]);
  assign t[67] = ~(t[126]);
  assign t[68] = ~(t[111]);
  assign t[69] = ~(t[127]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[90] & t[91]);
  assign t[72] = ~(t[129]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[92] & t[93]);
  assign t[75] = ~(t[94] & t[95]);
  assign t[76] = ~(t[96] & t[131]);
  assign t[77] = ~(t[122] & t[121]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[97] & t[98]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] & t[100]);
  assign t[85] = ~(t[101] & t[102]);
  assign t[86] = ~(t[103] & t[137]);
  assign t[87] = ~(t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[141]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[106] & t[107]);
  assign t[97] = ~(t[134] & t[133]);
  assign t[98] = ~(t[144]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[110];
endmodule

module R1ind192(x, y);
 input [94:0] x;
 output y;

 wire [152:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[100] = t[132] ^ x[40];
  assign t[101] = t[133] ^ x[45];
  assign t[102] = t[134] ^ x[47];
  assign t[103] = t[135] ^ x[51];
  assign t[104] = t[136] ^ x[54];
  assign t[105] = t[137] ^ x[56];
  assign t[106] = t[138] ^ x[59];
  assign t[107] = t[139] ^ x[61];
  assign t[108] = t[140] ^ x[66];
  assign t[109] = t[141] ^ x[68];
  assign t[10] = x[18] ^ x[19];
  assign t[110] = t[142] ^ x[72];
  assign t[111] = t[143] ^ x[75];
  assign t[112] = t[144] ^ x[77];
  assign t[113] = t[145] ^ x[79];
  assign t[114] = t[146] ^ x[81];
  assign t[115] = t[147] ^ x[83];
  assign t[116] = t[148] ^ x[85];
  assign t[117] = t[149] ^ x[88];
  assign t[118] = t[150] ^ x[90];
  assign t[119] = t[151] ^ x[92];
  assign t[11] = t[92] ? x[18] : x[19];
  assign t[120] = t[152] ^ x[94];
  assign t[121] = (x[0] & x[1]);
  assign t[122] = (x[6] & x[7]);
  assign t[123] = (x[9] & x[10]);
  assign t[124] = (x[12] & x[13]);
  assign t[125] = (x[15] & x[16]);
  assign t[126] = (x[20] & x[21]);
  assign t[127] = (x[20] & x[23]);
  assign t[128] = (x[27] & x[28]);
  assign t[129] = (x[27] & x[30]);
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = (x[20] & x[34]);
  assign t[131] = (x[36] & x[37]);
  assign t[132] = (x[36] & x[39]);
  assign t[133] = (x[43] & x[44]);
  assign t[134] = (x[43] & x[46]);
  assign t[135] = (x[27] & x[50]);
  assign t[136] = (x[52] & x[53]);
  assign t[137] = (x[52] & x[55]);
  assign t[138] = (x[57] & x[58]);
  assign t[139] = (x[57] & x[60]);
  assign t[13] = x[4] ? t[18] : t[17];
  assign t[140] = (x[64] & x[65]);
  assign t[141] = (x[64] & x[67]);
  assign t[142] = (x[36] & x[71]);
  assign t[143] = (x[73] & x[74]);
  assign t[144] = (x[73] & x[76]);
  assign t[145] = (x[43] & x[78]);
  assign t[146] = (x[52] & x[80]);
  assign t[147] = (x[57] & x[82]);
  assign t[148] = (x[64] & x[84]);
  assign t[149] = (x[86] & x[87]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (x[86] & x[89]);
  assign t[151] = (x[73] & x[91]);
  assign t[152] = (x[86] & x[93]);
  assign t[15] = x[4] ? t[22] : t[21];
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = t[27] ^ t[21];
  assign t[19] = x[4] ? t[29] : t[28];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = x[4] ? t[31] : t[30];
  assign t[21] = ~(t[32] & t[33]);
  assign t[22] = t[34] ^ t[35];
  assign t[23] = x[4] ? t[37] : t[36];
  assign t[24] = x[4] ? t[39] : t[38];
  assign t[25] = ~(t[94] & t[40]);
  assign t[26] = ~(t[95] & t[41]);
  assign t[27] = t[42] ? x[26] : x[25];
  assign t[28] = ~(t[43] & t[44]);
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[31] = t[49] ^ t[30];
  assign t[32] = ~(t[96] & t[50]);
  assign t[33] = ~(t[97] & t[51]);
  assign t[34] = t[42] ? x[33] : x[32];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[36];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = t[59] ^ t[60];
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[98]);
  assign t[41] = ~(t[98] & t[61]);
  assign t[42] = ~(t[62]);
  assign t[43] = ~(t[99] & t[63]);
  assign t[44] = ~(t[100] & t[64]);
  assign t[45] = t[42] ? x[42] : x[41];
  assign t[46] = ~(t[65] & t[66]);
  assign t[47] = ~(t[101] & t[67]);
  assign t[48] = ~(t[102] & t[68]);
  assign t[49] = t[42] ? x[49] : x[48];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = ~(t[103]);
  assign t[51] = ~(t[103] & t[69]);
  assign t[52] = ~(t[104] & t[70]);
  assign t[53] = ~(t[105] & t[71]);
  assign t[54] = ~(t[106] & t[72]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = t[92] ? x[63] : x[62];
  assign t[57] = ~(t[108] & t[74]);
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = t[92] ? x[70] : x[69];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = ~(t[76] & t[77]);
  assign t[61] = ~(t[94]);
  assign t[62] = ~(t[92]);
  assign t[63] = ~(t[110]);
  assign t[64] = ~(t[110] & t[78]);
  assign t[65] = ~(t[111] & t[79]);
  assign t[66] = ~(t[112] & t[80]);
  assign t[67] = ~(t[113]);
  assign t[68] = ~(t[113] & t[81]);
  assign t[69] = ~(t[96]);
  assign t[6] = ~(t[90] & t[91]);
  assign t[70] = ~(t[114]);
  assign t[71] = ~(t[114] & t[82]);
  assign t[72] = ~(t[115]);
  assign t[73] = ~(t[115] & t[83]);
  assign t[74] = ~(t[116]);
  assign t[75] = ~(t[116] & t[84]);
  assign t[76] = ~(t[117] & t[85]);
  assign t[77] = ~(t[118] & t[86]);
  assign t[78] = ~(t[99]);
  assign t[79] = ~(t[119]);
  assign t[7] = ~(t[92] & t[93]);
  assign t[80] = ~(t[119] & t[87]);
  assign t[81] = ~(t[101]);
  assign t[82] = ~(t[104]);
  assign t[83] = ~(t[106]);
  assign t[84] = ~(t[108]);
  assign t[85] = ~(t[120]);
  assign t[86] = ~(t[120] & t[88]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[117]);
  assign t[89] = t[121] ^ x[2];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[122] ^ x[8];
  assign t[91] = t[123] ^ x[11];
  assign t[92] = t[124] ^ x[14];
  assign t[93] = t[125] ^ x[17];
  assign t[94] = t[126] ^ x[22];
  assign t[95] = t[127] ^ x[24];
  assign t[96] = t[128] ^ x[29];
  assign t[97] = t[129] ^ x[31];
  assign t[98] = t[130] ^ x[35];
  assign t[99] = t[131] ^ x[38];
  assign t[9] = ~(t[13] ^ t[14]);
  assign y = t[0] ? t[1] : t[89];
endmodule

module R1ind193(x, y);
 input [112:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = ~(t[211] | t[212]);
  assign t[101] = ~(t[223]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[141] | t[142]);
  assign t[104] = ~(t[143] | t[144]);
  assign t[105] = ~(t[225]);
  assign t[106] = ~(t[226]);
  assign t[107] = ~(t[145] | t[146]);
  assign t[108] = ~(t[147] | t[148]);
  assign t[109] = ~(t[227] | t[149]);
  assign t[10] = ~(x[3]);
  assign t[110] = t[150] ? x[84] : x[83];
  assign t[111] = ~(t[151] & t[152]);
  assign t[112] = ~(t[228]);
  assign t[113] = ~(t[229]);
  assign t[114] = ~(t[153] | t[154]);
  assign t[115] = t[203] ? x[90] : x[89];
  assign t[116] = t[155] | t[156];
  assign t[117] = ~(t[203]);
  assign t[118] = ~(t[157] & t[204]);
  assign t[119] = ~(t[158] & t[159]);
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[120] = ~(t[76] | t[160]);
  assign t[121] = ~(t[76] | t[161]);
  assign t[122] = t[204] & t[162];
  assign t[123] = t[158] | t[157];
  assign t[124] = ~(t[163] & t[159]);
  assign t[125] = ~(x[4] & t[164]);
  assign t[126] = ~(t[158] & t[204]);
  assign t[127] = ~(t[157] & t[159]);
  assign t[128] = ~(t[203]);
  assign t[129] = ~(t[139]);
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[130] = ~(t[230]);
  assign t[131] = ~(t[217] | t[218]);
  assign t[132] = ~(t[165] | t[143]);
  assign t[133] = ~(t[166] | t[167]);
  assign t[134] = ~(t[231]);
  assign t[135] = ~(t[219] | t[220]);
  assign t[136] = ~(t[232]);
  assign t[137] = ~(t[233]);
  assign t[138] = ~(t[168] | t[169]);
  assign t[139] = ~(t[170] | t[143]);
  assign t[13] = x[4] ? t[22] : t[21];
  assign t[140] = ~(t[171] | t[172]);
  assign t[141] = ~(t[234]);
  assign t[142] = ~(t[223] | t[224]);
  assign t[143] = ~(t[117] | t[173]);
  assign t[144] = t[174] | t[175];
  assign t[145] = ~(t[235]);
  assign t[146] = ~(t[225] | t[226]);
  assign t[147] = ~(t[236]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[176] | t[177]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[150] = ~(t[128]);
  assign t[151] = ~(t[155] | t[178]);
  assign t[152] = ~(t[46]);
  assign t[153] = ~(t[238]);
  assign t[154] = ~(t[228] | t[229]);
  assign t[155] = ~(t[179] & t[180]);
  assign t[156] = ~(t[181] & t[85]);
  assign t[157] = x[4] & t[202];
  assign t[158] = ~(x[4] | t[202]);
  assign t[159] = ~(t[204]);
  assign t[15] = ~(t[201] & t[202]);
  assign t[160] = t[201] ? t[118] : t[119];
  assign t[161] = t[201] ? t[183] : t[182];
  assign t[162] = ~(t[117] | t[201]);
  assign t[163] = ~(x[4] | t[184]);
  assign t[164] = ~(t[202] | t[159]);
  assign t[165] = ~(t[117] | t[185]);
  assign t[166] = ~(t[30]);
  assign t[167] = ~(t[76] | t[186]);
  assign t[168] = ~(t[239]);
  assign t[169] = ~(t[232] | t[233]);
  assign t[16] = ~(t[203] & t[204]);
  assign t[170] = ~(t[117] | t[187]);
  assign t[171] = ~(t[188] & t[189]);
  assign t[172] = ~(t[79] & t[190]);
  assign t[173] = t[201] ? t[124] : t[183];
  assign t[174] = ~(t[76] | t[191]);
  assign t[175] = ~(t[179]);
  assign t[176] = ~(t[240]);
  assign t[177] = ~(t[236] | t[237]);
  assign t[178] = ~(t[192] & t[190]);
  assign t[179] = ~(t[162] & t[193]);
  assign t[17] = x[4] ? t[26] : t[25];
  assign t[180] = ~(t[164] & t[194]);
  assign t[181] = ~(t[46] | t[174]);
  assign t[182] = ~(t[204] & t[163]);
  assign t[183] = ~(x[4] & t[195]);
  assign t[184] = ~(t[202]);
  assign t[185] = t[201] ? t[119] : t[127];
  assign t[186] = t[201] ? t[182] : t[183];
  assign t[187] = t[201] ? t[127] : t[119];
  assign t[188] = ~(t[165] | t[196]);
  assign t[189] = ~(t[117] & t[197]);
  assign t[18] = ~(t[27] ^ t[28]);
  assign t[190] = t[117] | t[198];
  assign t[191] = t[201] ? t[126] : t[127];
  assign t[192] = ~(t[143]);
  assign t[193] = ~(t[182] & t[125]);
  assign t[194] = t[76] & t[201];
  assign t[195] = ~(t[202] | t[204]);
  assign t[196] = ~(t[76] | t[199]);
  assign t[197] = ~(t[183] & t[182]);
  assign t[198] = t[201] ? t[183] : t[124];
  assign t[199] = t[201] ? t[124] : t[125];
  assign t[19] = t[203] ? x[6] : x[7];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[200] = t[241] ^ x[2];
  assign t[201] = t[242] ^ x[10];
  assign t[202] = t[243] ^ x[13];
  assign t[203] = t[244] ^ x[16];
  assign t[204] = t[245] ^ x[19];
  assign t[205] = t[246] ^ x[22];
  assign t[206] = t[247] ^ x[25];
  assign t[207] = t[248] ^ x[27];
  assign t[208] = t[249] ^ x[29];
  assign t[209] = t[250] ^ x[34];
  assign t[20] = ~(t[29] & t[30]);
  assign t[210] = t[251] ^ x[37];
  assign t[211] = t[252] ^ x[39];
  assign t[212] = t[253] ^ x[41];
  assign t[213] = t[254] ^ x[44];
  assign t[214] = t[255] ^ x[49];
  assign t[215] = t[256] ^ x[52];
  assign t[216] = t[257] ^ x[54];
  assign t[217] = t[258] ^ x[56];
  assign t[218] = t[259] ^ x[58];
  assign t[219] = t[260] ^ x[62];
  assign t[21] = ~(t[31] | t[32]);
  assign t[220] = t[261] ^ x[64];
  assign t[221] = t[262] ^ x[67];
  assign t[222] = t[263] ^ x[71];
  assign t[223] = t[264] ^ x[73];
  assign t[224] = t[265] ^ x[75];
  assign t[225] = t[266] ^ x[77];
  assign t[226] = t[267] ^ x[79];
  assign t[227] = t[268] ^ x[82];
  assign t[228] = t[269] ^ x[86];
  assign t[229] = t[270] ^ x[88];
  assign t[22] = ~(t[25] ^ t[33]);
  assign t[230] = t[271] ^ x[92];
  assign t[231] = t[272] ^ x[94];
  assign t[232] = t[273] ^ x[96];
  assign t[233] = t[274] ^ x[98];
  assign t[234] = t[275] ^ x[100];
  assign t[235] = t[276] ^ x[102];
  assign t[236] = t[277] ^ x[104];
  assign t[237] = t[278] ^ x[106];
  assign t[238] = t[279] ^ x[108];
  assign t[239] = t[280] ^ x[110];
  assign t[23] = x[4] ? t[35] : t[34];
  assign t[240] = t[281] ^ x[112];
  assign t[241] = (x[0] & x[1]);
  assign t[242] = (x[8] & x[9]);
  assign t[243] = (x[11] & x[12]);
  assign t[244] = (x[14] & x[15]);
  assign t[245] = (x[17] & x[18]);
  assign t[246] = (x[20] & x[21]);
  assign t[247] = (x[23] & x[24]);
  assign t[248] = (x[20] & x[26]);
  assign t[249] = (x[20] & x[28]);
  assign t[24] = x[4] ? t[37] : t[36];
  assign t[250] = (x[32] & x[33]);
  assign t[251] = (x[35] & x[36]);
  assign t[252] = (x[23] & x[38]);
  assign t[253] = (x[23] & x[40]);
  assign t[254] = (x[42] & x[43]);
  assign t[255] = (x[47] & x[48]);
  assign t[256] = (x[50] & x[51]);
  assign t[257] = (x[20] & x[53]);
  assign t[258] = (x[32] & x[55]);
  assign t[259] = (x[32] & x[57]);
  assign t[25] = ~(t[38] | t[39]);
  assign t[260] = (x[35] & x[61]);
  assign t[261] = (x[35] & x[63]);
  assign t[262] = (x[65] & x[66]);
  assign t[263] = (x[23] & x[70]);
  assign t[264] = (x[42] & x[72]);
  assign t[265] = (x[42] & x[74]);
  assign t[266] = (x[47] & x[76]);
  assign t[267] = (x[47] & x[78]);
  assign t[268] = (x[80] & x[81]);
  assign t[269] = (x[50] & x[85]);
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = (x[50] & x[87]);
  assign t[271] = (x[32] & x[91]);
  assign t[272] = (x[35] & x[93]);
  assign t[273] = (x[65] & x[95]);
  assign t[274] = (x[65] & x[97]);
  assign t[275] = (x[42] & x[99]);
  assign t[276] = (x[47] & x[101]);
  assign t[277] = (x[80] & x[103]);
  assign t[278] = (x[80] & x[105]);
  assign t[279] = (x[50] & x[107]);
  assign t[27] = x[4] ? t[43] : t[42];
  assign t[280] = (x[65] & x[109]);
  assign t[281] = (x[80] & x[111]);
  assign t[28] = x[4] ? t[45] : t[44];
  assign t[29] = ~(t[46] | t[47]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[32] = ~(t[205] | t[52]);
  assign t[33] = ~(t[53] ^ t[54]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[35] = ~(t[34] ^ t[57]);
  assign t[36] = ~(t[58] | t[59]);
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[39] = ~(t[206] | t[64]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[65] | t[66]);
  assign t[41] = ~(t[67] ^ t[68]);
  assign t[42] = ~(t[69] | t[70]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[45] = ~(t[44] ^ t[75]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[47] = ~(t[78] & t[79]);
  assign t[48] = ~(t[76] | t[80]);
  assign t[49] = ~(t[76] | t[81]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[207]);
  assign t[51] = ~(t[208]);
  assign t[52] = ~(t[82] | t[83]);
  assign t[53] = t[84] ? x[31] : x[30];
  assign t[54] = ~(t[85] & t[86]);
  assign t[55] = ~(t[87] | t[88]);
  assign t[56] = ~(t[209] | t[89]);
  assign t[57] = ~(t[90] ^ t[91]);
  assign t[58] = ~(t[92] | t[93]);
  assign t[59] = ~(t[210] | t[94]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[97] ^ t[98]);
  assign t[62] = ~(t[211]);
  assign t[63] = ~(t[212]);
  assign t[64] = ~(t[99] | t[100]);
  assign t[65] = ~(t[101] | t[102]);
  assign t[66] = ~(t[213] | t[103]);
  assign t[67] = t[203] ? x[46] : x[45];
  assign t[68] = ~(t[29] & t[104]);
  assign t[69] = ~(t[105] | t[106]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = ~(t[214] | t[107]);
  assign t[71] = ~(t[108] | t[109]);
  assign t[72] = ~(t[110] ^ t[111]);
  assign t[73] = ~(t[112] | t[113]);
  assign t[74] = ~(t[215] | t[114]);
  assign t[75] = ~(t[115] ^ t[116]);
  assign t[76] = ~(t[117]);
  assign t[77] = t[201] ? t[119] : t[118];
  assign t[78] = ~(t[120] | t[121]);
  assign t[79] = ~(t[122] & t[123]);
  assign t[7] = ~(t[13] ^ t[14]);
  assign t[80] = t[201] ? t[125] : t[124];
  assign t[81] = t[201] ? t[127] : t[126];
  assign t[82] = ~(t[216]);
  assign t[83] = ~(t[207] | t[208]);
  assign t[84] = ~(t[128]);
  assign t[85] = ~(t[121] | t[49]);
  assign t[86] = ~(t[122] | t[129]);
  assign t[87] = ~(t[217]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[130] | t[131]);
  assign t[8] = x[6] ^ x[7];
  assign t[90] = t[84] ? x[60] : x[59];
  assign t[91] = ~(t[132] & t[133]);
  assign t[92] = ~(t[219]);
  assign t[93] = ~(t[220]);
  assign t[94] = ~(t[134] | t[135]);
  assign t[95] = ~(t[136] | t[137]);
  assign t[96] = ~(t[221] | t[138]);
  assign t[97] = t[84] ? x[69] : x[68];
  assign t[98] = ~(t[139] & t[140]);
  assign t[99] = ~(t[222]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = t[0] ? t[1] : t[200];
endmodule

module R1ind194(x, y);
 input [12:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[10] ^ t[1];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = (x[1] & x[2]);
  assign t[15] = (x[4] & x[5]);
  assign t[16] = (x[7] & x[8]);
  assign t[17] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[11]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[3] = ~(t[12]);
  assign t[4] = ~(t[5] & t[13]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[11] & t[10]);
  assign t[9] = ~(t[13] & t[12]);
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind195(x, y);
 input [12:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[9] ^ t[1]);
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[9];
  assign t[12] = t[16] ^ x[12];
  assign t[13] = (x[1] & x[2]);
  assign t[14] = (x[4] & x[5]);
  assign t[15] = (x[7] & x[8]);
  assign t[16] = (x[10] & x[11]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[10]);
  assign t[3] = ~(t[4] & t[11]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(x[0]);
  assign t[7] = ~(t[9] & t[12]);
  assign t[8] = ~(t[11] & t[10]);
  assign t[9] = t[13] ^ x[3];
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind196(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = t[7] ^ t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = ~(t[8] & t[7]);
  assign t[7] = t[11] ^ x[3];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[9];
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind197(x, y);
 input [12:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[6] ^ t[1]);
  assign t[10] = (x[1] & x[2]);
  assign t[11] = (x[4] & x[5]);
  assign t[12] = (x[7] & x[8]);
  assign t[13] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(x[0]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[6] & t[9]);
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[6];
  assign t[8] = t[12] ^ x[9];
  assign t[9] = t[13] ^ x[12];
  assign y = ~(x[0] | t[0]);
endmodule

module R1_ind(x, y);
 input [496:0] x;
 output [197:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[7], x[6], x[3]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[9], x[8], x[3]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[11], x[10], x[3]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[14], x[13], x[12]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[16], x[15], x[12]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[18], x[17], x[12]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[20], x[19], x[12]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[23], x[22], x[21]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[25], x[24], x[21]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[27], x[26], x[21]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[29], x[28], x[21]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[32], x[31], x[30]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[34], x[33], x[30]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[36], x[35], x[30]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[38], x[37], x[30]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[41], x[40], x[39]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[43], x[42], x[39]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[45], x[44], x[39]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[47], x[46], x[39]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[50], x[49], x[48]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[52], x[51], x[48]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[54], x[53], x[48]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[56], x[55], x[48]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[59], x[58], x[57]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[61], x[60], x[57]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[63], x[62], x[57]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[65], x[64], x[57]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[68], x[67], x[66]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[70], x[69], x[66]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[72], x[71], x[66]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[74], x[73], x[66]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[77], x[76], x[75]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[79], x[78], x[75]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[81], x[80], x[75]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[83], x[82], x[75]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[86], x[85], x[84]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[88], x[87], x[84]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[90], x[89], x[84]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[92], x[91], x[84]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[95], x[94], x[93]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[97], x[96], x[93]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[99], x[98], x[93]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[101], x[100], x[93]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[104], x[103], x[102]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[106], x[105], x[102]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[108], x[107], x[102]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[110], x[109], x[102]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[113], x[112], x[111]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[115], x[114], x[111]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[117], x[116], x[111]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[119], x[118], x[111]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[122], x[121], x[120]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[124], x[123], x[120]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[126], x[125], x[120]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[128], x[127], x[120]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[131], x[130], x[129]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[133], x[132], x[129]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[135], x[134], x[129]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[137], x[136], x[129]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[140], x[139], x[138]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[142], x[141], x[138]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[144], x[143], x[138]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[146], x[145], x[138]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[159], x[158]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[153], x[152], x[155], x[154], x[157], x[156], x[149], x[161], x[160]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[155], x[154], x[153], x[152], x[157], x[156], x[151], x[150], x[149], x[163], x[162]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[167], x[166], x[176], x[175]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[170], x[169], x[172], x[171], x[174], x[173], x[166], x[178], x[177]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[172], x[171], x[170], x[169], x[174], x[173], x[168], x[167], x[166], x[180], x[179]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[193], x[192]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[187], x[186], x[189], x[188], x[191], x[190], x[183], x[195], x[194]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[189], x[188], x[187], x[186], x[191], x[190], x[185], x[184], x[183], x[197], x[196]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[210], x[209]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[204], x[203], x[206], x[205], x[208], x[207], x[200], x[212], x[211]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[206], x[205], x[204], x[203], x[208], x[207], x[202], x[201], x[200], x[214], x[213]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[227], x[226]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[221], x[220], x[223], x[222], x[225], x[224], x[217], x[229], x[228]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[223], x[222], x[221], x[220], x[225], x[224], x[219], x[218], x[217], x[231], x[230]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[244], x[243]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[238], x[237], x[240], x[239], x[242], x[241], x[234], x[246], x[245]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[240], x[239], x[238], x[237], x[242], x[241], x[236], x[235], x[234], x[248], x[247]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[259], x[258], x[257], x[256], x[255], x[254], x[253], x[252], x[251], x[261], x[260]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[255], x[254], x[257], x[256], x[259], x[258], x[251], x[263], x[262]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[257], x[256], x[255], x[254], x[259], x[258], x[253], x[252], x[251], x[265], x[264]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[278], x[277]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[272], x[271], x[274], x[273], x[276], x[275], x[268], x[280], x[279]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[274], x[273], x[272], x[271], x[276], x[275], x[270], x[269], x[268], x[282], x[281]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[293], x[292], x[291], x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[283]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[293], x[292], x[291], x[290], x[289], x[288], x[287], x[286], x[285], x[295], x[294]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[289], x[288], x[291], x[290], x[293], x[292], x[285], x[297], x[296]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[291], x[290], x[289], x[288], x[293], x[292], x[287], x[286], x[285], x[299], x[298]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[300]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[310], x[309], x[308], x[307], x[306], x[305], x[304], x[303], x[302], x[312], x[311]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[306], x[305], x[308], x[307], x[310], x[309], x[302], x[314], x[313]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[308], x[307], x[306], x[305], x[310], x[309], x[304], x[303], x[302], x[316], x[315]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[327], x[326], x[325], x[324], x[323], x[322], x[321], x[320], x[319], x[318], x[317]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[327], x[326], x[325], x[324], x[323], x[322], x[321], x[320], x[319], x[329], x[328]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[323], x[322], x[325], x[324], x[327], x[326], x[319], x[331], x[330]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[325], x[324], x[323], x[322], x[327], x[326], x[321], x[320], x[319], x[333], x[332]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[336], x[335], x[334]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[337], x[336], x[346], x[345]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[340], x[339], x[342], x[341], x[344], x[343], x[336], x[348], x[347]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[342], x[341], x[340], x[339], x[344], x[343], x[338], x[337], x[336], x[350], x[349]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[352], x[351]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[363], x[362]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[357], x[356], x[359], x[358], x[361], x[360], x[353], x[365], x[364]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[359], x[358], x[357], x[356], x[361], x[360], x[355], x[354], x[353], x[367], x[366]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[378], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[370], x[369], x[368]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[378], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[370], x[380], x[379]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[374], x[373], x[376], x[375], x[378], x[377], x[370], x[382], x[381]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[376], x[375], x[374], x[373], x[378], x[377], x[372], x[371], x[370], x[384], x[383]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[388], x[387], x[386], x[385]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[388], x[387], x[397], x[396]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[391], x[390], x[393], x[392], x[395], x[394], x[387], x[399], x[398]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[393], x[392], x[391], x[390], x[395], x[394], x[389], x[388], x[387], x[401], x[400]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[405], x[404], x[403], x[402]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[405], x[404], x[414], x[413]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[408], x[407], x[410], x[409], x[412], x[411], x[404], x[416], x[415]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[410], x[409], x[408], x[407], x[412], x[411], x[406], x[405], x[404], x[418], x[417]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[191], x[190], x[208], x[207], x[189], x[188], x[187], x[186], x[242], x[241], x[206], x[205], x[204], x[203], x[412], x[411], x[174], x[173], x[185], x[184], x[183], x[240], x[239], x[238], x[237], x[202], x[201], x[200], x[410], x[409], x[408], x[407], x[172], x[171], x[170], x[169], x[327], x[326], x[182], x[181], x[236], x[235], x[234], x[199], x[198], x[406], x[405], x[404], x[168], x[167], x[166], x[325], x[324], x[323], x[322], x[165], x[164], x[321], x[320], x[319], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[148], x[147], x[433], x[432], x[431], x[153], x[152], x[149]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[191], x[190], x[208], x[207], x[189], x[188], x[187], x[186], x[242], x[241], x[206], x[205], x[204], x[203], x[412], x[411], x[174], x[173], x[185], x[184], x[183], x[240], x[239], x[238], x[237], x[202], x[201], x[200], x[410], x[409], x[408], x[407], x[172], x[171], x[170], x[169], x[327], x[326], x[193], x[192], x[236], x[235], x[234], x[210], x[209], x[406], x[405], x[404], x[168], x[167], x[166], x[325], x[324], x[323], x[322], x[176], x[175], x[321], x[320], x[319], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[159], x[158], x[434], x[432], x[431], x[157], x[156], x[149]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[187], x[186], x[204], x[203], x[189], x[188], x[191], x[190], x[183], x[238], x[237], x[206], x[205], x[208], x[207], x[200], x[408], x[407], x[170], x[169], x[195], x[194], x[240], x[239], x[242], x[241], x[234], x[212], x[211], x[410], x[409], x[412], x[411], x[404], x[172], x[171], x[174], x[173], x[166], x[323], x[322], x[178], x[177], x[325], x[324], x[327], x[326], x[319], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[161], x[160], x[435], x[432], x[431], x[151], x[150], x[149]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[206], x[205], x[189], x[188], x[204], x[203], x[208], x[207], x[410], x[409], x[187], x[186], x[191], x[190], x[240], x[239], x[172], x[171], x[214], x[213], x[202], x[201], x[200], x[408], x[407], x[412], x[411], x[197], x[196], x[185], x[184], x[183], x[238], x[237], x[242], x[241], x[170], x[169], x[174], x[173], x[325], x[324], x[406], x[405], x[404], x[236], x[235], x[234], x[180], x[179], x[168], x[167], x[166], x[323], x[322], x[327], x[326], x[321], x[320], x[319], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[163], x[162], x[436], x[432], x[431], x[155], x[154], x[149]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[191], x[190], x[208], x[207], x[189], x[188], x[187], x[186], x[242], x[241], x[206], x[205], x[204], x[203], x[412], x[411], x[225], x[224], x[395], x[394], x[259], x[258], x[185], x[184], x[183], x[240], x[239], x[238], x[237], x[202], x[201], x[200], x[410], x[409], x[408], x[407], x[157], x[156], x[223], x[222], x[221], x[220], x[393], x[392], x[391], x[390], x[257], x[256], x[255], x[254], x[344], x[343], x[182], x[181], x[236], x[235], x[234], x[199], x[198], x[406], x[405], x[404], x[155], x[154], x[153], x[152], x[233], x[232], x[219], x[218], x[217], x[216], x[215], x[389], x[388], x[387], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[148], x[147], x[151], x[150], x[149], x[250], x[249], x[338], x[337], x[336], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[165], x[164], x[437], x[432], x[431], x[170], x[169], x[166]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[191], x[190], x[208], x[207], x[189], x[188], x[187], x[186], x[242], x[241], x[206], x[205], x[204], x[203], x[412], x[411], x[225], x[224], x[395], x[394], x[259], x[258], x[185], x[184], x[183], x[240], x[239], x[238], x[237], x[202], x[201], x[200], x[410], x[409], x[408], x[407], x[157], x[156], x[223], x[222], x[221], x[220], x[393], x[392], x[391], x[390], x[257], x[256], x[255], x[254], x[344], x[343], x[193], x[192], x[236], x[235], x[234], x[210], x[209], x[406], x[405], x[404], x[155], x[154], x[153], x[152], x[244], x[243], x[219], x[218], x[217], x[227], x[226], x[389], x[388], x[387], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[159], x[158], x[151], x[150], x[149], x[261], x[260], x[338], x[337], x[336], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[176], x[175], x[438], x[432], x[431], x[174], x[173], x[166]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[187], x[186], x[204], x[203], x[189], x[188], x[191], x[190], x[183], x[238], x[237], x[206], x[205], x[208], x[207], x[200], x[408], x[407], x[391], x[390], x[221], x[220], x[255], x[254], x[195], x[194], x[240], x[239], x[242], x[241], x[234], x[212], x[211], x[410], x[409], x[412], x[411], x[404], x[153], x[152], x[229], x[228], x[393], x[392], x[395], x[394], x[387], x[246], x[245], x[223], x[222], x[225], x[224], x[217], x[257], x[256], x[259], x[258], x[251], x[340], x[339], x[161], x[160], x[155], x[154], x[157], x[156], x[149], x[263], x[262], x[342], x[341], x[344], x[343], x[336], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[178], x[177], x[439], x[432], x[431], x[168], x[167], x[166]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[206], x[205], x[189], x[188], x[204], x[203], x[208], x[207], x[410], x[409], x[187], x[186], x[191], x[190], x[240], x[239], x[223], x[222], x[393], x[392], x[257], x[256], x[214], x[213], x[202], x[201], x[200], x[408], x[407], x[412], x[411], x[197], x[196], x[185], x[184], x[183], x[238], x[237], x[242], x[241], x[155], x[154], x[248], x[247], x[221], x[220], x[225], x[224], x[231], x[230], x[391], x[390], x[395], x[394], x[255], x[254], x[259], x[258], x[342], x[341], x[406], x[405], x[404], x[236], x[235], x[234], x[163], x[162], x[153], x[152], x[157], x[156], x[219], x[218], x[217], x[389], x[388], x[387], x[265], x[264], x[253], x[252], x[251], x[340], x[339], x[344], x[343], x[151], x[150], x[149], x[338], x[337], x[336], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[180], x[179], x[440], x[432], x[431], x[172], x[171], x[166]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[174], x[173], x[361], x[360], x[172], x[171], x[170], x[169], x[327], x[326], x[157], x[156], x[208], x[207], x[378], x[377], x[359], x[358], x[357], x[356], x[276], x[275], x[168], x[167], x[166], x[325], x[324], x[323], x[322], x[155], x[154], x[153], x[152], x[206], x[205], x[204], x[203], x[412], x[411], x[376], x[375], x[374], x[373], x[355], x[354], x[353], x[274], x[273], x[272], x[271], x[293], x[292], x[165], x[164], x[321], x[320], x[319], x[148], x[147], x[151], x[150], x[149], x[202], x[201], x[200], x[410], x[409], x[408], x[407], x[368], x[369], x[372], x[371], x[370], x[351], x[352], x[270], x[269], x[268], x[291], x[290], x[289], x[288], x[199], x[198], x[406], x[405], x[404], x[402], x[403], x[287], x[286], x[285], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[182], x[181], x[441], x[432], x[431], x[187], x[186], x[183]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[174], x[173], x[361], x[360], x[172], x[171], x[170], x[169], x[327], x[326], x[157], x[156], x[208], x[207], x[378], x[377], x[359], x[358], x[357], x[356], x[276], x[275], x[168], x[167], x[166], x[325], x[324], x[323], x[322], x[155], x[154], x[153], x[152], x[206], x[205], x[204], x[203], x[412], x[411], x[376], x[375], x[374], x[373], x[355], x[354], x[353], x[274], x[273], x[272], x[271], x[293], x[292], x[176], x[175], x[321], x[320], x[319], x[159], x[158], x[151], x[150], x[149], x[202], x[201], x[200], x[410], x[409], x[408], x[407], x[379], x[380], x[372], x[371], x[370], x[362], x[363], x[270], x[269], x[268], x[291], x[290], x[289], x[288], x[210], x[209], x[406], x[405], x[404], x[413], x[414], x[287], x[286], x[285], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[193], x[192], x[442], x[432], x[431], x[191], x[190], x[183]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[170], x[169], x[357], x[356], x[153], x[152], x[172], x[171], x[174], x[173], x[166], x[323], x[322], x[204], x[203], x[359], x[358], x[361], x[360], x[353], x[272], x[271], x[374], x[373], x[161], x[160], x[155], x[154], x[157], x[156], x[149], x[178], x[177], x[325], x[324], x[327], x[326], x[319], x[206], x[205], x[208], x[207], x[200], x[408], x[407], x[364], x[365], x[274], x[273], x[276], x[275], x[268], x[382], x[381], x[376], x[375], x[378], x[377], x[370], x[289], x[288], x[212], x[211], x[410], x[409], x[412], x[411], x[404], x[415], x[416], x[291], x[290], x[293], x[292], x[285], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[195], x[194], x[443], x[432], x[431], x[185], x[184], x[183]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[172], x[171], x[359], x[358], x[170], x[169], x[174], x[173], x[325], x[324], x[155], x[154], x[206], x[205], x[376], x[375], x[357], x[356], x[361], x[360], x[274], x[273], x[180], x[179], x[168], x[167], x[166], x[323], x[322], x[327], x[326], x[163], x[162], x[153], x[152], x[157], x[156], x[204], x[203], x[208], x[207], x[410], x[409], x[384], x[383], x[374], x[373], x[378], x[377], x[366], x[367], x[355], x[354], x[353], x[272], x[271], x[276], x[275], x[291], x[290], x[321], x[320], x[319], x[151], x[150], x[149], x[214], x[213], x[202], x[201], x[200], x[408], x[407], x[412], x[411], x[372], x[371], x[370], x[270], x[269], x[268], x[417], x[418], x[289], x[288], x[293], x[292], x[406], x[405], x[404], x[287], x[286], x[285], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[197], x[196], x[444], x[432], x[431], x[189], x[188], x[183]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[174], x[173], x[344], x[343], x[172], x[171], x[170], x[169], x[327], x[326], x[157], x[156], x[191], x[190], x[361], x[360], x[342], x[341], x[340], x[339], x[259], x[258], x[293], x[292], x[168], x[167], x[166], x[325], x[324], x[323], x[322], x[155], x[154], x[153], x[152], x[189], x[188], x[187], x[186], x[242], x[241], x[359], x[358], x[357], x[356], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[291], x[290], x[289], x[288], x[310], x[309], x[165], x[164], x[321], x[320], x[319], x[148], x[147], x[151], x[150], x[149], x[185], x[184], x[183], x[240], x[239], x[238], x[237], x[317], x[318], x[355], x[354], x[353], x[334], x[335], x[253], x[252], x[251], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[182], x[181], x[236], x[235], x[234], x[283], x[284], x[304], x[303], x[302], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[199], x[198], x[445], x[432], x[431], x[204], x[203], x[200]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[174], x[173], x[344], x[343], x[172], x[171], x[170], x[169], x[327], x[326], x[157], x[156], x[191], x[190], x[361], x[360], x[342], x[341], x[340], x[339], x[259], x[258], x[293], x[292], x[168], x[167], x[166], x[325], x[324], x[323], x[322], x[155], x[154], x[153], x[152], x[189], x[188], x[187], x[186], x[242], x[241], x[359], x[358], x[357], x[356], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[291], x[290], x[289], x[288], x[310], x[309], x[176], x[175], x[321], x[320], x[319], x[159], x[158], x[151], x[150], x[149], x[185], x[184], x[183], x[240], x[239], x[238], x[237], x[328], x[329], x[355], x[354], x[353], x[345], x[346], x[253], x[252], x[251], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[193], x[192], x[236], x[235], x[234], x[294], x[295], x[304], x[303], x[302], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[210], x[209], x[446], x[432], x[431], x[208], x[207], x[200]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[170], x[169], x[340], x[339], x[153], x[152], x[172], x[171], x[174], x[173], x[166], x[323], x[322], x[187], x[186], x[357], x[356], x[342], x[341], x[344], x[343], x[336], x[255], x[254], x[289], x[288], x[161], x[160], x[155], x[154], x[157], x[156], x[149], x[178], x[177], x[325], x[324], x[327], x[326], x[319], x[189], x[188], x[191], x[190], x[183], x[238], x[237], x[330], x[331], x[359], x[358], x[361], x[360], x[353], x[347], x[348], x[257], x[256], x[259], x[258], x[251], x[291], x[290], x[293], x[292], x[285], x[306], x[305], x[195], x[194], x[240], x[239], x[242], x[241], x[234], x[296], x[297], x[308], x[307], x[310], x[309], x[302], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[212], x[211], x[447], x[432], x[431], x[202], x[201], x[200]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[172], x[171], x[342], x[341], x[170], x[169], x[174], x[173], x[325], x[324], x[155], x[154], x[189], x[188], x[340], x[339], x[344], x[343], x[257], x[256], x[359], x[358], x[291], x[290], x[180], x[179], x[168], x[167], x[166], x[323], x[322], x[327], x[326], x[163], x[162], x[153], x[152], x[157], x[156], x[187], x[186], x[191], x[190], x[240], x[239], x[349], x[350], x[338], x[337], x[336], x[255], x[254], x[259], x[258], x[332], x[333], x[357], x[356], x[361], x[360], x[289], x[288], x[293], x[292], x[308], x[307], x[321], x[320], x[319], x[151], x[150], x[149], x[197], x[196], x[185], x[184], x[183], x[238], x[237], x[242], x[241], x[253], x[252], x[251], x[355], x[354], x[353], x[298], x[299], x[287], x[286], x[285], x[306], x[305], x[310], x[309], x[236], x[235], x[234], x[304], x[303], x[302], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[214], x[213], x[448], x[432], x[431], x[206], x[205], x[200]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[259], x[258], x[276], x[275], x[242], x[241], x[257], x[256], x[255], x[254], x[344], x[343], x[274], x[273], x[272], x[271], x[174], x[173], x[240], x[239], x[238], x[237], x[225], x[224], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[270], x[269], x[268], x[172], x[171], x[170], x[169], x[395], x[394], x[236], x[235], x[234], x[223], x[222], x[250], x[249], x[338], x[337], x[336], x[266], x[267], x[168], x[167], x[166], x[393], x[392], x[391], x[390], x[233], x[232], x[219], x[218], x[389], x[388], x[387], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[216], x[215], x[449], x[432], x[431], x[221], x[220], x[217]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[259], x[258], x[276], x[275], x[242], x[241], x[257], x[256], x[255], x[254], x[344], x[343], x[274], x[273], x[272], x[271], x[174], x[173], x[240], x[239], x[238], x[237], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[270], x[269], x[268], x[172], x[171], x[170], x[169], x[395], x[394], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[261], x[260], x[338], x[337], x[336], x[277], x[278], x[168], x[167], x[166], x[393], x[392], x[391], x[390], x[244], x[243], x[219], x[218], x[389], x[388], x[387], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[227], x[226], x[450], x[432], x[431], x[225], x[224], x[217]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[255], x[254], x[272], x[271], x[238], x[237], x[257], x[256], x[259], x[258], x[251], x[340], x[339], x[274], x[273], x[276], x[275], x[268], x[170], x[169], x[240], x[239], x[242], x[241], x[234], x[221], x[220], x[263], x[262], x[342], x[341], x[344], x[343], x[336], x[279], x[280], x[172], x[171], x[174], x[173], x[166], x[391], x[390], x[246], x[245], x[223], x[222], x[225], x[224], x[393], x[392], x[395], x[394], x[387], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[229], x[228], x[451], x[432], x[431], x[219], x[218], x[217]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[274], x[273], x[257], x[256], x[240], x[239], x[272], x[271], x[276], x[275], x[172], x[171], x[255], x[254], x[259], x[258], x[342], x[341], x[238], x[237], x[242], x[241], x[281], x[282], x[270], x[269], x[268], x[170], x[169], x[174], x[173], x[265], x[264], x[253], x[252], x[251], x[340], x[339], x[344], x[343], x[393], x[392], x[248], x[247], x[236], x[235], x[234], x[221], x[220], x[225], x[224], x[168], x[167], x[166], x[338], x[337], x[336], x[391], x[390], x[395], x[394], x[219], x[218], x[389], x[388], x[387], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[231], x[230], x[452], x[432], x[431], x[223], x[222], x[217]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[259], x[258], x[276], x[275], x[257], x[256], x[255], x[254], x[344], x[343], x[274], x[273], x[272], x[271], x[174], x[173], x[225], x[224], x[327], x[326], x[157], x[156], x[208], x[207], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[270], x[269], x[268], x[172], x[171], x[170], x[169], x[223], x[222], x[221], x[220], x[395], x[394], x[325], x[324], x[323], x[322], x[155], x[154], x[153], x[152], x[206], x[205], x[204], x[203], x[412], x[411], x[250], x[249], x[338], x[337], x[336], x[266], x[267], x[168], x[167], x[166], x[219], x[218], x[217], x[393], x[392], x[391], x[390], x[165], x[164], x[321], x[320], x[319], x[148], x[147], x[151], x[150], x[149], x[202], x[201], x[200], x[410], x[409], x[408], x[407], x[216], x[215], x[389], x[388], x[387], x[199], x[198], x[406], x[405], x[404], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[233], x[232], x[453], x[432], x[431], x[238], x[237], x[234]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[259], x[258], x[276], x[275], x[257], x[256], x[255], x[254], x[344], x[343], x[274], x[273], x[272], x[271], x[174], x[173], x[225], x[224], x[327], x[326], x[157], x[156], x[208], x[207], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[270], x[269], x[268], x[172], x[171], x[170], x[169], x[223], x[222], x[221], x[220], x[395], x[394], x[325], x[324], x[323], x[322], x[155], x[154], x[153], x[152], x[206], x[205], x[204], x[203], x[412], x[411], x[261], x[260], x[338], x[337], x[336], x[277], x[278], x[168], x[167], x[166], x[219], x[218], x[217], x[393], x[392], x[391], x[390], x[176], x[175], x[321], x[320], x[319], x[159], x[158], x[151], x[150], x[149], x[202], x[201], x[200], x[410], x[409], x[408], x[407], x[227], x[226], x[389], x[388], x[387], x[210], x[209], x[406], x[405], x[404], x[244], x[243], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[454], x[432], x[431], x[242], x[241], x[234]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[255], x[254], x[272], x[271], x[257], x[256], x[259], x[258], x[251], x[340], x[339], x[274], x[273], x[276], x[275], x[268], x[170], x[169], x[221], x[220], x[153], x[152], x[323], x[322], x[204], x[203], x[263], x[262], x[342], x[341], x[344], x[343], x[336], x[279], x[280], x[172], x[171], x[174], x[173], x[166], x[223], x[222], x[225], x[224], x[217], x[391], x[390], x[161], x[160], x[155], x[154], x[157], x[156], x[149], x[178], x[177], x[325], x[324], x[327], x[326], x[319], x[206], x[205], x[208], x[207], x[200], x[408], x[407], x[229], x[228], x[393], x[392], x[395], x[394], x[387], x[212], x[211], x[410], x[409], x[412], x[411], x[404], x[246], x[245], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[455], x[432], x[431], x[236], x[235], x[234]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[274], x[273], x[257], x[256], x[272], x[271], x[276], x[275], x[172], x[171], x[255], x[254], x[259], x[258], x[342], x[341], x[223], x[222], x[325], x[324], x[155], x[154], x[206], x[205], x[281], x[282], x[270], x[269], x[268], x[170], x[169], x[174], x[173], x[265], x[264], x[253], x[252], x[251], x[340], x[339], x[344], x[343], x[221], x[220], x[225], x[224], x[393], x[392], x[180], x[179], x[323], x[322], x[327], x[326], x[163], x[162], x[153], x[152], x[157], x[156], x[204], x[203], x[208], x[207], x[410], x[409], x[168], x[167], x[166], x[338], x[337], x[336], x[231], x[230], x[219], x[218], x[217], x[391], x[390], x[395], x[394], x[321], x[320], x[319], x[151], x[150], x[149], x[214], x[213], x[202], x[201], x[200], x[408], x[407], x[412], x[411], x[389], x[388], x[387], x[406], x[405], x[404], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[248], x[247], x[456], x[432], x[431], x[240], x[239], x[234]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[242], x[241], x[293], x[292], x[240], x[239], x[238], x[237], x[225], x[224], x[395], x[394], x[276], x[275], x[208], x[207], x[291], x[290], x[289], x[288], x[310], x[309], x[327], x[326], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[393], x[392], x[391], x[390], x[274], x[273], x[272], x[271], x[174], x[173], x[206], x[205], x[204], x[203], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[325], x[324], x[323], x[322], x[361], x[360], x[233], x[232], x[219], x[218], x[217], x[216], x[215], x[389], x[388], x[387], x[270], x[269], x[268], x[172], x[171], x[170], x[169], x[300], x[301], x[202], x[201], x[200], x[283], x[284], x[304], x[303], x[302], x[321], x[320], x[319], x[359], x[358], x[357], x[356], x[266], x[267], x[168], x[167], x[166], x[317], x[318], x[355], x[354], x[353], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[250], x[249], x[457], x[432], x[431], x[255], x[254], x[251]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[242], x[241], x[293], x[292], x[240], x[239], x[238], x[237], x[225], x[224], x[395], x[394], x[276], x[275], x[208], x[207], x[291], x[290], x[289], x[288], x[310], x[309], x[327], x[326], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[393], x[392], x[391], x[390], x[274], x[273], x[272], x[271], x[174], x[173], x[206], x[205], x[204], x[203], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[325], x[324], x[323], x[322], x[361], x[360], x[244], x[243], x[219], x[218], x[217], x[227], x[226], x[389], x[388], x[387], x[270], x[269], x[268], x[172], x[171], x[170], x[169], x[311], x[312], x[202], x[201], x[200], x[294], x[295], x[304], x[303], x[302], x[321], x[320], x[319], x[359], x[358], x[357], x[356], x[277], x[278], x[168], x[167], x[166], x[328], x[329], x[355], x[354], x[353], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[261], x[260], x[458], x[432], x[431], x[259], x[258], x[251]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[238], x[237], x[289], x[288], x[391], x[390], x[240], x[239], x[242], x[241], x[234], x[221], x[220], x[272], x[271], x[291], x[290], x[293], x[292], x[285], x[306], x[305], x[204], x[203], x[323], x[322], x[229], x[228], x[393], x[392], x[395], x[394], x[387], x[246], x[245], x[223], x[222], x[225], x[224], x[217], x[274], x[273], x[276], x[275], x[268], x[170], x[169], x[296], x[297], x[308], x[307], x[310], x[309], x[302], x[313], x[314], x[206], x[205], x[208], x[207], x[200], x[325], x[324], x[327], x[326], x[319], x[357], x[356], x[279], x[280], x[172], x[171], x[174], x[173], x[166], x[330], x[331], x[359], x[358], x[361], x[360], x[353], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[263], x[262], x[459], x[432], x[431], x[253], x[252], x[251]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[240], x[239], x[291], x[290], x[238], x[237], x[242], x[241], x[223], x[222], x[393], x[392], x[274], x[273], x[206], x[205], x[289], x[288], x[293], x[292], x[308], x[307], x[325], x[324], x[248], x[247], x[236], x[235], x[234], x[221], x[220], x[225], x[224], x[231], x[230], x[391], x[390], x[395], x[394], x[272], x[271], x[276], x[275], x[172], x[171], x[315], x[316], x[204], x[203], x[208], x[207], x[298], x[299], x[287], x[286], x[285], x[306], x[305], x[310], x[309], x[323], x[322], x[327], x[326], x[359], x[358], x[219], x[218], x[217], x[389], x[388], x[387], x[281], x[282], x[270], x[269], x[268], x[170], x[169], x[174], x[173], x[202], x[201], x[200], x[304], x[303], x[302], x[332], x[333], x[321], x[320], x[319], x[357], x[356], x[361], x[360], x[168], x[167], x[166], x[355], x[354], x[353], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[265], x[264], x[460], x[432], x[431], x[257], x[256], x[251]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[242], x[241], x[412], x[411], x[240], x[239], x[238], x[237], x[225], x[224], x[395], x[394], x[259], x[258], x[191], x[190], x[410], x[409], x[408], x[407], x[293], x[292], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[393], x[392], x[391], x[390], x[257], x[256], x[255], x[254], x[344], x[343], x[189], x[188], x[187], x[186], x[406], x[405], x[404], x[291], x[290], x[289], x[288], x[378], x[377], x[233], x[232], x[219], x[218], x[217], x[216], x[215], x[389], x[388], x[387], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[386], x[385], x[185], x[184], x[183], x[402], x[403], x[287], x[286], x[285], x[376], x[375], x[374], x[373], x[250], x[249], x[338], x[337], x[336], x[368], x[369], x[372], x[371], x[370], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[267], x[266], x[461], x[432], x[431], x[272], x[271], x[268]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[242], x[241], x[412], x[411], x[240], x[239], x[238], x[237], x[225], x[224], x[395], x[394], x[259], x[258], x[191], x[190], x[410], x[409], x[408], x[407], x[293], x[292], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[393], x[392], x[391], x[390], x[257], x[256], x[255], x[254], x[344], x[343], x[189], x[188], x[187], x[186], x[406], x[405], x[404], x[291], x[290], x[289], x[288], x[378], x[377], x[244], x[243], x[219], x[218], x[217], x[227], x[226], x[389], x[388], x[387], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[396], x[397], x[185], x[184], x[183], x[413], x[414], x[287], x[286], x[285], x[376], x[375], x[374], x[373], x[261], x[260], x[338], x[337], x[336], x[379], x[380], x[372], x[371], x[370], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[278], x[277], x[462], x[432], x[431], x[276], x[275], x[268]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[238], x[237], x[408], x[407], x[391], x[390], x[240], x[239], x[242], x[241], x[234], x[221], x[220], x[255], x[254], x[187], x[186], x[410], x[409], x[412], x[411], x[404], x[289], x[288], x[229], x[228], x[393], x[392], x[395], x[394], x[387], x[246], x[245], x[223], x[222], x[225], x[224], x[217], x[257], x[256], x[259], x[258], x[251], x[340], x[339], x[398], x[399], x[189], x[188], x[191], x[190], x[183], x[415], x[416], x[291], x[290], x[293], x[292], x[285], x[374], x[373], x[263], x[262], x[342], x[341], x[344], x[343], x[336], x[382], x[381], x[376], x[375], x[378], x[377], x[370], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[280], x[279], x[463], x[432], x[431], x[270], x[269], x[268]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[240], x[239], x[410], x[409], x[238], x[237], x[242], x[241], x[223], x[222], x[393], x[392], x[257], x[256], x[408], x[407], x[412], x[411], x[291], x[290], x[189], x[188], x[248], x[247], x[236], x[235], x[234], x[221], x[220], x[225], x[224], x[231], x[230], x[391], x[390], x[395], x[394], x[255], x[254], x[259], x[258], x[342], x[341], x[417], x[418], x[406], x[405], x[404], x[289], x[288], x[293], x[292], x[400], x[401], x[187], x[186], x[191], x[190], x[376], x[375], x[219], x[218], x[217], x[389], x[388], x[387], x[265], x[264], x[253], x[252], x[251], x[340], x[339], x[344], x[343], x[287], x[286], x[285], x[185], x[184], x[183], x[384], x[383], x[374], x[373], x[378], x[377], x[338], x[337], x[336], x[372], x[371], x[370], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[282], x[281], x[464], x[432], x[431], x[274], x[273], x[268]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[327], x[326], x[344], x[343], x[325], x[324], x[323], x[322], x[361], x[360], x[342], x[341], x[340], x[339], x[259], x[258], x[310], x[309], x[378], x[377], x[276], x[275], x[395], x[394], x[321], x[320], x[319], x[359], x[358], x[357], x[356], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[308], x[307], x[306], x[305], x[208], x[207], x[376], x[375], x[374], x[373], x[274], x[273], x[272], x[271], x[393], x[392], x[391], x[390], x[191], x[190], x[317], x[318], x[355], x[354], x[353], x[334], x[335], x[253], x[252], x[251], x[304], x[303], x[302], x[206], x[205], x[204], x[203], x[368], x[369], x[372], x[371], x[370], x[351], x[352], x[270], x[269], x[268], x[389], x[388], x[387], x[189], x[188], x[187], x[186], x[300], x[301], x[202], x[201], x[200], x[386], x[385], x[185], x[184], x[183], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[284], x[283], x[465], x[432], x[431], x[289], x[288], x[285]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[327], x[326], x[344], x[343], x[325], x[324], x[323], x[322], x[361], x[360], x[342], x[341], x[340], x[339], x[259], x[258], x[310], x[309], x[378], x[377], x[276], x[275], x[395], x[394], x[321], x[320], x[319], x[359], x[358], x[357], x[356], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[308], x[307], x[306], x[305], x[208], x[207], x[376], x[375], x[374], x[373], x[274], x[273], x[272], x[271], x[393], x[392], x[391], x[390], x[191], x[190], x[328], x[329], x[355], x[354], x[353], x[345], x[346], x[253], x[252], x[251], x[304], x[303], x[302], x[206], x[205], x[204], x[203], x[379], x[380], x[372], x[371], x[370], x[362], x[363], x[270], x[269], x[268], x[389], x[388], x[387], x[189], x[188], x[187], x[186], x[311], x[312], x[202], x[201], x[200], x[396], x[397], x[185], x[184], x[183], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[295], x[294], x[466], x[432], x[431], x[293], x[292], x[285]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[323], x[322], x[340], x[339], x[325], x[324], x[327], x[326], x[319], x[357], x[356], x[342], x[341], x[344], x[343], x[336], x[255], x[254], x[306], x[305], x[272], x[271], x[374], x[373], x[391], x[390], x[330], x[331], x[359], x[358], x[361], x[360], x[353], x[347], x[348], x[257], x[256], x[259], x[258], x[251], x[308], x[307], x[310], x[309], x[302], x[204], x[203], x[364], x[365], x[274], x[273], x[276], x[275], x[268], x[382], x[381], x[376], x[375], x[378], x[377], x[370], x[393], x[392], x[395], x[394], x[387], x[187], x[186], x[313], x[314], x[206], x[205], x[208], x[207], x[200], x[398], x[399], x[189], x[188], x[191], x[190], x[183], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[297], x[296], x[467], x[432], x[431], x[287], x[286], x[285]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[342], x[341], x[325], x[324], x[340], x[339], x[344], x[343], x[257], x[256], x[323], x[322], x[327], x[326], x[359], x[358], x[308], x[307], x[376], x[375], x[274], x[273], x[393], x[392], x[349], x[350], x[338], x[337], x[336], x[255], x[254], x[259], x[258], x[332], x[333], x[321], x[320], x[319], x[357], x[356], x[361], x[360], x[306], x[305], x[310], x[309], x[206], x[205], x[384], x[383], x[374], x[373], x[378], x[377], x[366], x[367], x[272], x[271], x[276], x[275], x[391], x[390], x[395], x[394], x[189], x[188], x[253], x[252], x[251], x[355], x[354], x[353], x[315], x[316], x[304], x[303], x[302], x[204], x[203], x[208], x[207], x[372], x[371], x[370], x[270], x[269], x[268], x[400], x[401], x[389], x[388], x[387], x[187], x[186], x[191], x[190], x[202], x[201], x[200], x[185], x[184], x[183], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[299], x[298], x[468], x[432], x[431], x[291], x[290], x[285]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[327], x[326], x[344], x[343], x[293], x[292], x[325], x[324], x[323], x[322], x[361], x[360], x[342], x[341], x[340], x[339], x[259], x[258], x[291], x[290], x[289], x[288], x[310], x[309], x[321], x[320], x[319], x[359], x[358], x[357], x[356], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[208], x[207], x[287], x[286], x[285], x[308], x[307], x[317], x[318], x[355], x[354], x[353], x[334], x[335], x[253], x[252], x[251], x[206], x[205], x[204], x[203], x[283], x[284], x[304], x[303], x[202], x[201], x[200], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[301], x[300], x[469], x[432], x[431], x[306], x[305], x[302]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[327], x[326], x[344], x[343], x[293], x[292], x[325], x[324], x[323], x[322], x[361], x[360], x[342], x[341], x[340], x[339], x[259], x[258], x[291], x[290], x[289], x[288], x[321], x[320], x[319], x[359], x[358], x[357], x[356], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[208], x[207], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[328], x[329], x[355], x[354], x[353], x[345], x[346], x[253], x[252], x[251], x[206], x[205], x[204], x[203], x[294], x[295], x[304], x[303], x[202], x[201], x[200], x[430], x[429], x[428], x[424], x[423], x[422], x[421], x[420], x[419], x[427], x[426], x[425], x[312], x[311], x[470], x[432], x[431], x[310], x[309], x[302]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[323], x[322], x[340], x[339], x[289], x[288], x[325], x[324], x[327], x[326], x[319], x[357], x[356], x[342], x[341], x[344], x[343], x[336], x[255], x[254], x[291], x[290], x[293], x[292], x[285], x[306], x[305], x[330], x[331], x[359], x[358], x[361], x[360], x[353], x[347], x[348], x[257], x[256], x[259], x[258], x[251], x[204], x[203], x[296], x[297], x[308], x[307], x[310], x[309], x[206], x[205], x[208], x[207], x[200], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[314], x[313], x[471], x[432], x[431], x[304], x[303], x[302]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[342], x[341], x[325], x[324], x[291], x[290], x[340], x[339], x[344], x[343], x[257], x[256], x[323], x[322], x[327], x[326], x[359], x[358], x[289], x[288], x[293], x[292], x[349], x[350], x[338], x[337], x[336], x[255], x[254], x[259], x[258], x[332], x[333], x[321], x[320], x[319], x[357], x[356], x[361], x[360], x[206], x[205], x[298], x[299], x[287], x[286], x[285], x[306], x[305], x[310], x[309], x[253], x[252], x[251], x[355], x[354], x[353], x[204], x[203], x[208], x[207], x[304], x[303], x[202], x[201], x[200], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[316], x[315], x[472], x[432], x[431], x[308], x[307], x[302]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[293], x[292], x[191], x[190], x[208], x[207], x[291], x[290], x[289], x[288], x[310], x[309], x[344], x[343], x[189], x[188], x[187], x[186], x[242], x[241], x[412], x[411], x[206], x[205], x[204], x[203], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[342], x[341], x[340], x[339], x[259], x[258], x[185], x[184], x[183], x[240], x[239], x[238], x[237], x[410], x[409], x[408], x[407], x[157], x[156], x[300], x[301], x[202], x[201], x[200], x[283], x[284], x[304], x[303], x[302], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[182], x[181], x[236], x[235], x[234], x[199], x[198], x[406], x[405], x[404], x[155], x[154], x[153], x[152], x[334], x[335], x[253], x[252], x[251], x[148], x[147], x[151], x[150], x[149], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[318], x[317], x[473], x[432], x[431], x[323], x[322], x[319]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[293], x[292], x[191], x[190], x[208], x[207], x[291], x[290], x[289], x[288], x[310], x[309], x[344], x[343], x[189], x[188], x[187], x[186], x[242], x[241], x[412], x[411], x[206], x[205], x[204], x[203], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[342], x[341], x[340], x[339], x[259], x[258], x[185], x[184], x[183], x[240], x[239], x[238], x[237], x[410], x[409], x[408], x[407], x[157], x[156], x[311], x[312], x[202], x[201], x[200], x[294], x[295], x[304], x[303], x[302], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[193], x[192], x[236], x[235], x[234], x[210], x[209], x[406], x[405], x[404], x[155], x[154], x[153], x[152], x[345], x[346], x[253], x[252], x[251], x[159], x[158], x[151], x[150], x[149], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[329], x[328], x[474], x[432], x[431], x[327], x[326], x[319]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[289], x[288], x[187], x[186], x[291], x[290], x[293], x[292], x[285], x[306], x[305], x[204], x[203], x[340], x[339], x[189], x[188], x[191], x[190], x[183], x[238], x[237], x[408], x[407], x[296], x[297], x[308], x[307], x[310], x[309], x[302], x[313], x[314], x[206], x[205], x[208], x[207], x[200], x[342], x[341], x[344], x[343], x[336], x[255], x[254], x[195], x[194], x[240], x[239], x[242], x[241], x[234], x[212], x[211], x[410], x[409], x[412], x[411], x[404], x[153], x[152], x[347], x[348], x[257], x[256], x[259], x[258], x[251], x[161], x[160], x[155], x[154], x[157], x[156], x[149], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[331], x[330], x[475], x[432], x[431], x[321], x[320], x[319]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[291], x[290], x[189], x[188], x[206], x[205], x[289], x[288], x[293], x[292], x[308], x[307], x[342], x[341], x[410], x[409], x[187], x[186], x[191], x[190], x[240], x[239], x[315], x[316], x[204], x[203], x[208], x[207], x[298], x[299], x[287], x[286], x[285], x[306], x[305], x[310], x[309], x[340], x[339], x[344], x[343], x[257], x[256], x[214], x[213], x[408], x[407], x[412], x[411], x[197], x[196], x[185], x[184], x[183], x[238], x[237], x[242], x[241], x[155], x[154], x[202], x[201], x[200], x[304], x[303], x[302], x[349], x[350], x[338], x[337], x[336], x[255], x[254], x[259], x[258], x[406], x[405], x[404], x[236], x[235], x[234], x[163], x[162], x[153], x[152], x[157], x[156], x[253], x[252], x[251], x[151], x[150], x[149], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[333], x[332], x[476], x[432], x[431], x[325], x[324], x[319]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[293], x[292], x[242], x[241], x[208], x[207], x[291], x[290], x[289], x[288], x[310], x[309], x[327], x[326], x[240], x[239], x[238], x[237], x[225], x[224], x[395], x[394], x[276], x[275], x[206], x[205], x[204], x[203], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[325], x[324], x[323], x[322], x[361], x[360], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[393], x[392], x[391], x[390], x[274], x[273], x[272], x[271], x[174], x[173], x[300], x[301], x[202], x[201], x[200], x[283], x[284], x[304], x[303], x[302], x[321], x[320], x[319], x[359], x[358], x[357], x[356], x[233], x[232], x[219], x[218], x[217], x[216], x[215], x[389], x[388], x[387], x[270], x[269], x[268], x[172], x[171], x[170], x[169], x[317], x[318], x[355], x[354], x[353], x[266], x[267], x[168], x[167], x[166], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[335], x[334], x[477], x[432], x[431], x[340], x[339], x[336]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[293], x[292], x[242], x[241], x[208], x[207], x[291], x[290], x[289], x[288], x[310], x[309], x[327], x[326], x[240], x[239], x[238], x[237], x[225], x[224], x[395], x[394], x[276], x[275], x[206], x[205], x[204], x[203], x[287], x[286], x[285], x[308], x[307], x[306], x[305], x[325], x[324], x[323], x[322], x[361], x[360], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[393], x[392], x[391], x[390], x[274], x[273], x[272], x[271], x[174], x[173], x[311], x[312], x[202], x[201], x[200], x[294], x[295], x[304], x[303], x[302], x[321], x[320], x[319], x[359], x[358], x[357], x[356], x[244], x[243], x[219], x[218], x[217], x[227], x[226], x[389], x[388], x[387], x[270], x[269], x[268], x[172], x[171], x[170], x[169], x[328], x[329], x[355], x[354], x[353], x[277], x[278], x[168], x[167], x[166], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[346], x[345], x[478], x[432], x[431], x[344], x[343], x[336]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[289], x[288], x[238], x[237], x[291], x[290], x[293], x[292], x[285], x[306], x[305], x[204], x[203], x[323], x[322], x[391], x[390], x[240], x[239], x[242], x[241], x[234], x[221], x[220], x[272], x[271], x[296], x[297], x[308], x[307], x[310], x[309], x[302], x[313], x[314], x[206], x[205], x[208], x[207], x[200], x[325], x[324], x[327], x[326], x[319], x[357], x[356], x[229], x[228], x[393], x[392], x[395], x[394], x[387], x[246], x[245], x[223], x[222], x[225], x[224], x[217], x[274], x[273], x[276], x[275], x[268], x[170], x[169], x[330], x[331], x[359], x[358], x[361], x[360], x[353], x[279], x[280], x[172], x[171], x[174], x[173], x[166], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[348], x[347], x[479], x[432], x[431], x[338], x[337], x[336]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[291], x[290], x[240], x[239], x[206], x[205], x[289], x[288], x[293], x[292], x[308], x[307], x[325], x[324], x[238], x[237], x[242], x[241], x[223], x[222], x[393], x[392], x[274], x[273], x[315], x[316], x[204], x[203], x[208], x[207], x[298], x[299], x[287], x[286], x[285], x[306], x[305], x[310], x[309], x[323], x[322], x[327], x[326], x[359], x[358], x[248], x[247], x[236], x[235], x[234], x[221], x[220], x[225], x[224], x[231], x[230], x[391], x[390], x[395], x[394], x[272], x[271], x[276], x[275], x[172], x[171], x[202], x[201], x[200], x[304], x[303], x[302], x[332], x[333], x[321], x[320], x[319], x[357], x[356], x[361], x[360], x[219], x[218], x[217], x[389], x[388], x[387], x[281], x[282], x[270], x[269], x[268], x[170], x[169], x[174], x[173], x[355], x[354], x[353], x[168], x[167], x[166], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[350], x[349], x[480], x[432], x[431], x[342], x[341], x[336]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[395], x[394], x[412], x[411], x[393], x[392], x[391], x[390], x[191], x[190], x[410], x[409], x[408], x[407], x[293], x[292], x[208], x[207], x[310], x[309], x[344], x[343], x[389], x[388], x[387], x[189], x[188], x[187], x[186], x[406], x[405], x[404], x[291], x[290], x[289], x[288], x[378], x[377], x[206], x[205], x[204], x[203], x[308], x[307], x[306], x[305], x[342], x[341], x[340], x[339], x[259], x[258], x[386], x[385], x[185], x[184], x[183], x[402], x[403], x[287], x[286], x[285], x[376], x[375], x[374], x[373], x[300], x[301], x[202], x[201], x[200], x[283], x[284], x[304], x[303], x[302], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[368], x[369], x[372], x[371], x[370], x[334], x[335], x[253], x[252], x[251], x[352], x[351], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[481], x[432], x[431], x[357], x[356], x[353]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[395], x[394], x[412], x[411], x[393], x[392], x[391], x[390], x[191], x[190], x[410], x[409], x[408], x[407], x[293], x[292], x[208], x[207], x[310], x[309], x[344], x[343], x[389], x[388], x[387], x[189], x[188], x[187], x[186], x[406], x[405], x[404], x[291], x[290], x[289], x[288], x[378], x[377], x[206], x[205], x[204], x[203], x[308], x[307], x[306], x[305], x[342], x[341], x[340], x[339], x[259], x[258], x[396], x[397], x[185], x[184], x[183], x[413], x[414], x[287], x[286], x[285], x[376], x[375], x[374], x[373], x[311], x[312], x[202], x[201], x[200], x[294], x[295], x[304], x[303], x[302], x[338], x[337], x[336], x[257], x[256], x[255], x[254], x[379], x[380], x[372], x[371], x[370], x[345], x[346], x[253], x[252], x[251], x[363], x[362], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[482], x[432], x[431], x[361], x[360], x[353]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[391], x[390], x[408], x[407], x[393], x[392], x[395], x[394], x[387], x[187], x[186], x[410], x[409], x[412], x[411], x[404], x[289], x[288], x[306], x[305], x[204], x[203], x[340], x[339], x[398], x[399], x[189], x[188], x[191], x[190], x[183], x[415], x[416], x[291], x[290], x[293], x[292], x[285], x[374], x[373], x[296], x[297], x[308], x[307], x[310], x[309], x[302], x[313], x[314], x[206], x[205], x[208], x[207], x[200], x[342], x[341], x[344], x[343], x[336], x[255], x[254], x[382], x[381], x[376], x[375], x[378], x[377], x[370], x[347], x[348], x[257], x[256], x[259], x[258], x[251], x[365], x[364], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[483], x[432], x[431], x[355], x[354], x[353]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[410], x[409], x[393], x[392], x[408], x[407], x[412], x[411], x[291], x[290], x[391], x[390], x[395], x[394], x[189], x[188], x[206], x[205], x[308], x[307], x[342], x[341], x[417], x[418], x[406], x[405], x[404], x[289], x[288], x[293], x[292], x[400], x[401], x[389], x[388], x[387], x[187], x[186], x[191], x[190], x[376], x[375], x[315], x[316], x[204], x[203], x[208], x[207], x[298], x[299], x[306], x[305], x[310], x[309], x[340], x[339], x[344], x[343], x[257], x[256], x[287], x[286], x[285], x[185], x[184], x[183], x[384], x[383], x[374], x[373], x[378], x[377], x[202], x[201], x[200], x[304], x[303], x[302], x[349], x[350], x[338], x[337], x[336], x[255], x[254], x[259], x[258], x[372], x[371], x[370], x[253], x[252], x[251], x[367], x[366], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[484], x[432], x[431], x[359], x[358], x[353]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[395], x[394], x[412], x[411], x[393], x[392], x[391], x[390], x[191], x[190], x[410], x[409], x[408], x[407], x[293], x[292], x[361], x[360], x[389], x[388], x[387], x[189], x[188], x[187], x[186], x[406], x[405], x[404], x[291], x[290], x[289], x[288], x[359], x[358], x[357], x[356], x[276], x[275], x[386], x[385], x[185], x[184], x[183], x[402], x[403], x[287], x[286], x[285], x[355], x[354], x[353], x[274], x[273], x[272], x[271], x[351], x[352], x[270], x[269], x[268], x[369], x[368], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[485], x[432], x[431], x[374], x[373], x[370]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[395], x[394], x[412], x[411], x[393], x[392], x[391], x[390], x[191], x[190], x[410], x[409], x[408], x[407], x[293], x[292], x[361], x[360], x[389], x[388], x[387], x[189], x[188], x[187], x[186], x[406], x[405], x[404], x[291], x[290], x[289], x[288], x[359], x[358], x[357], x[356], x[276], x[275], x[396], x[397], x[185], x[184], x[183], x[413], x[414], x[287], x[286], x[285], x[355], x[354], x[353], x[274], x[273], x[272], x[271], x[362], x[363], x[270], x[269], x[268], x[380], x[379], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[486], x[432], x[431], x[378], x[377], x[370]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[391], x[390], x[408], x[407], x[393], x[392], x[395], x[394], x[387], x[187], x[186], x[410], x[409], x[412], x[411], x[404], x[289], x[288], x[357], x[356], x[398], x[399], x[189], x[188], x[191], x[190], x[183], x[415], x[416], x[291], x[290], x[293], x[292], x[285], x[359], x[358], x[361], x[360], x[353], x[272], x[271], x[364], x[365], x[274], x[273], x[276], x[275], x[268], x[382], x[381], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[487], x[432], x[431], x[372], x[371], x[370]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[410], x[409], x[393], x[392], x[408], x[407], x[412], x[411], x[291], x[290], x[391], x[390], x[395], x[394], x[189], x[188], x[359], x[358], x[417], x[418], x[406], x[405], x[404], x[289], x[288], x[293], x[292], x[400], x[401], x[389], x[388], x[387], x[187], x[186], x[191], x[190], x[357], x[356], x[361], x[360], x[274], x[273], x[287], x[286], x[285], x[185], x[184], x[183], x[366], x[367], x[355], x[354], x[353], x[272], x[271], x[276], x[275], x[270], x[269], x[268], x[384], x[383], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[488], x[432], x[431], x[376], x[375], x[370]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[361], x[360], x[259], x[258], x[378], x[377], x[359], x[358], x[357], x[356], x[276], x[275], x[412], x[411], x[257], x[256], x[255], x[254], x[344], x[343], x[174], x[173], x[242], x[241], x[376], x[375], x[374], x[373], x[355], x[354], x[353], x[274], x[273], x[272], x[271], x[410], x[409], x[408], x[407], x[293], x[292], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[172], x[171], x[170], x[169], x[240], x[239], x[238], x[237], x[225], x[224], x[368], x[369], x[372], x[371], x[370], x[351], x[352], x[270], x[269], x[268], x[406], x[405], x[404], x[291], x[290], x[289], x[288], x[250], x[249], x[338], x[337], x[336], x[266], x[267], x[168], x[167], x[166], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[402], x[403], x[287], x[286], x[285], x[233], x[232], x[219], x[218], x[217], x[386], x[385], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[489], x[432], x[431], x[391], x[390], x[387]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[361], x[360], x[259], x[258], x[378], x[377], x[359], x[358], x[357], x[356], x[276], x[275], x[412], x[411], x[257], x[256], x[255], x[254], x[344], x[343], x[174], x[173], x[242], x[241], x[376], x[375], x[374], x[373], x[355], x[354], x[353], x[274], x[273], x[272], x[271], x[410], x[409], x[408], x[407], x[293], x[292], x[253], x[252], x[251], x[342], x[341], x[340], x[339], x[172], x[171], x[170], x[169], x[240], x[239], x[238], x[237], x[225], x[224], x[379], x[380], x[372], x[371], x[370], x[362], x[363], x[270], x[269], x[268], x[406], x[405], x[404], x[291], x[290], x[289], x[288], x[261], x[260], x[338], x[337], x[336], x[277], x[278], x[168], x[167], x[166], x[236], x[235], x[234], x[223], x[222], x[221], x[220], x[413], x[414], x[287], x[286], x[285], x[244], x[243], x[219], x[218], x[217], x[397], x[396], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[490], x[432], x[431], x[395], x[394], x[387]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[357], x[356], x[255], x[254], x[359], x[358], x[361], x[360], x[353], x[272], x[271], x[374], x[373], x[408], x[407], x[257], x[256], x[259], x[258], x[251], x[340], x[339], x[170], x[169], x[238], x[237], x[364], x[365], x[274], x[273], x[276], x[275], x[268], x[382], x[381], x[376], x[375], x[378], x[377], x[370], x[410], x[409], x[412], x[411], x[404], x[289], x[288], x[263], x[262], x[342], x[341], x[344], x[343], x[336], x[279], x[280], x[172], x[171], x[174], x[173], x[166], x[240], x[239], x[242], x[241], x[234], x[221], x[220], x[415], x[416], x[291], x[290], x[293], x[292], x[285], x[246], x[245], x[223], x[222], x[225], x[224], x[217], x[399], x[398], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[491], x[432], x[431], x[389], x[388], x[387]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[359], x[358], x[257], x[256], x[376], x[375], x[357], x[356], x[361], x[360], x[274], x[273], x[410], x[409], x[172], x[171], x[255], x[254], x[259], x[258], x[342], x[341], x[240], x[239], x[384], x[383], x[374], x[373], x[378], x[377], x[366], x[367], x[355], x[354], x[353], x[272], x[271], x[276], x[275], x[408], x[407], x[412], x[411], x[291], x[290], x[281], x[282], x[170], x[169], x[174], x[173], x[265], x[264], x[253], x[252], x[251], x[340], x[339], x[344], x[343], x[238], x[237], x[242], x[241], x[223], x[222], x[372], x[371], x[370], x[270], x[269], x[268], x[417], x[418], x[406], x[405], x[404], x[289], x[288], x[293], x[292], x[168], x[167], x[166], x[338], x[337], x[336], x[248], x[247], x[236], x[235], x[234], x[221], x[220], x[225], x[224], x[287], x[286], x[285], x[219], x[218], x[217], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[401], x[400], x[492], x[432], x[431], x[393], x[392], x[387]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[361], x[360], x[174], x[173], x[378], x[377], x[359], x[358], x[357], x[356], x[276], x[275], x[395], x[394], x[172], x[171], x[170], x[169], x[327], x[326], x[157], x[156], x[376], x[375], x[374], x[373], x[355], x[354], x[353], x[274], x[273], x[272], x[271], x[393], x[392], x[391], x[390], x[191], x[190], x[168], x[167], x[166], x[325], x[324], x[323], x[322], x[155], x[154], x[153], x[152], x[242], x[241], x[368], x[369], x[372], x[371], x[370], x[351], x[352], x[270], x[269], x[268], x[389], x[388], x[387], x[189], x[188], x[187], x[186], x[165], x[164], x[321], x[320], x[319], x[148], x[147], x[151], x[150], x[149], x[240], x[239], x[238], x[237], x[386], x[385], x[185], x[184], x[183], x[182], x[181], x[236], x[235], x[234], x[403], x[402], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[493], x[432], x[431], x[408], x[407], x[404]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[361], x[360], x[174], x[173], x[378], x[377], x[359], x[358], x[357], x[356], x[276], x[275], x[395], x[394], x[172], x[171], x[170], x[169], x[327], x[326], x[157], x[156], x[376], x[375], x[374], x[373], x[355], x[354], x[353], x[274], x[273], x[272], x[271], x[393], x[392], x[391], x[390], x[191], x[190], x[168], x[167], x[166], x[325], x[324], x[323], x[322], x[155], x[154], x[153], x[152], x[242], x[241], x[379], x[380], x[372], x[371], x[370], x[362], x[363], x[270], x[269], x[268], x[389], x[388], x[387], x[189], x[188], x[187], x[186], x[176], x[175], x[321], x[320], x[319], x[159], x[158], x[151], x[150], x[149], x[240], x[239], x[238], x[237], x[396], x[397], x[185], x[184], x[183], x[193], x[192], x[236], x[235], x[234], x[430], x[429], x[428], x[424], x[423], x[422], x[421], x[420], x[419], x[427], x[426], x[425], x[414], x[413], x[494], x[432], x[431], x[412], x[411], x[404]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[357], x[356], x[170], x[169], x[359], x[358], x[361], x[360], x[353], x[272], x[271], x[374], x[373], x[391], x[390], x[153], x[152], x[172], x[171], x[174], x[173], x[166], x[323], x[322], x[364], x[365], x[274], x[273], x[276], x[275], x[268], x[382], x[381], x[376], x[375], x[378], x[377], x[370], x[393], x[392], x[395], x[394], x[387], x[187], x[186], x[161], x[160], x[155], x[154], x[157], x[156], x[149], x[178], x[177], x[325], x[324], x[327], x[326], x[319], x[238], x[237], x[398], x[399], x[189], x[188], x[191], x[190], x[183], x[195], x[194], x[240], x[239], x[242], x[241], x[234], x[416], x[415], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[495], x[432], x[431], x[406], x[405], x[404]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[359], x[358], x[172], x[171], x[376], x[375], x[357], x[356], x[361], x[360], x[274], x[273], x[393], x[392], x[170], x[169], x[174], x[173], x[325], x[324], x[155], x[154], x[384], x[383], x[374], x[373], x[378], x[377], x[366], x[367], x[355], x[354], x[353], x[272], x[271], x[276], x[275], x[391], x[390], x[395], x[394], x[189], x[188], x[180], x[179], x[168], x[167], x[166], x[323], x[322], x[327], x[326], x[163], x[162], x[153], x[152], x[157], x[156], x[240], x[239], x[372], x[371], x[370], x[270], x[269], x[268], x[400], x[401], x[389], x[388], x[387], x[187], x[186], x[191], x[190], x[321], x[320], x[319], x[151], x[150], x[149], x[197], x[196], x[238], x[237], x[242], x[241], x[185], x[184], x[183], x[236], x[235], x[234], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[418], x[417], x[496], x[432], x[431], x[410], x[409], x[404]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[427], x[426], x[425], x[430], x[429], x[428], x[421], x[420], x[419], x[424], x[423], x[422], x[431]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[424], x[423], x[422], x[427], x[426], x[425], x[430], x[429], x[428], x[421], x[420], x[419], x[431]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[424], x[423], x[422], x[421], x[420], x[419], x[427], x[426], x[425], x[430], x[429], x[428], x[431]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[430], x[429], x[428], x[424], x[423], x[422], x[421], x[420], x[419], x[427], x[426], x[425], x[431]}), .y(y[197]));
endmodule

module R2ind0(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[10] = (1'b0);
  assign t[11] = (x[0]);
  assign t[1] = (t[2] & ~t[3] & ~t[4] & ~t[5] & ~t[6]);
  assign t[2] = t[7] ^ x[5];
  assign t[3] = t[8] ^ x[1];
  assign t[4] = t[9] ^ x[2];
  assign t[5] = t[10] ^ x[3];
  assign t[6] = t[11] ^ x[4];
  assign t[7] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (1'b0);
  assign t[9] = (1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [11:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[14] ^ x[11];
  assign t[11] = (~t[15] & t[16]);
  assign t[12] = (~t[17] & t[18]);
  assign t[13] = (~t[19] & t[20]);
  assign t[14] = (~t[21] & t[22]);
  assign t[15] = t[23] ^ x[1];
  assign t[16] = t[24] ^ x[2];
  assign t[17] = t[25] ^ x[4];
  assign t[18] = t[26] ^ x[5];
  assign t[19] = t[27] ^ x[7];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[28] ^ x[8];
  assign t[21] = t[29] ^ x[10];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[24] = (x[0]);
  assign t[25] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[26] = (x[3]);
  assign t[27] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[6]);
  assign t[29] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (x[9]);
  assign t[3] = (t[7]);
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind6(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind7(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind8(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind9(x, y);
 input [11:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[14] ^ x[11];
  assign t[11] = (~t[15] & t[16]);
  assign t[12] = (~t[17] & t[18]);
  assign t[13] = (~t[19] & t[20]);
  assign t[14] = (~t[21] & t[22]);
  assign t[15] = t[23] ^ x[1];
  assign t[16] = t[24] ^ x[2];
  assign t[17] = t[25] ^ x[4];
  assign t[18] = t[26] ^ x[5];
  assign t[19] = t[27] ^ x[7];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[28] ^ x[8];
  assign t[21] = t[29] ^ x[10];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[24] = (x[0]);
  assign t[25] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[26] = (x[3]);
  assign t[27] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[6]);
  assign t[29] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (x[9]);
  assign t[3] = (t[7]);
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [12:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = ~(t[14] & t[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[3];
  assign t[16] = t[20] ^ x[6];
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[12];
  assign t[19] = (~t[23] & t[24]);
  assign t[1] = t[11] ^ t[2];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[3];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[6];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[3] & t[12]);
  assign t[30] = t[38] ^ x[12];
  assign t[31] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[1]);
  assign t[33] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[4]);
  assign t[35] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[7]);
  assign t[37] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[13]);
  assign t[5] = ~(t[6] & t[14]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(x[0]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind14(x, y);
 input [12:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = ~(t[14] & t[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[3];
  assign t[16] = t[20] ^ x[6];
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[12];
  assign t[19] = (~t[23] & t[24]);
  assign t[1] = t[11] ^ t[2];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[3];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[6];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[3] & t[12]);
  assign t[30] = t[38] ^ x[12];
  assign t[31] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[1]);
  assign t[33] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[4]);
  assign t[35] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[7]);
  assign t[37] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[13]);
  assign t[5] = ~(t[6] & t[14]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(x[0]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [12:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[3];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[12];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = ~(t[10] ^ t[2]);
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[1]);
  assign t[32] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[4]);
  assign t[34] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[7]);
  assign t[36] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[10]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[5] & t[12]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[10] & t[13]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind16(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind17(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind19(x, y);
 input [12:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[3];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[12];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = ~(t[10] ^ t[2]);
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[1]);
  assign t[32] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[4]);
  assign t[34] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[7]);
  assign t[36] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[10]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[5] & t[12]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[10] & t[13]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [12:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[3];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[9];
  assign t[15] = t[19] ^ x[12];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[8] ^ t[2];
  assign t[20] = t[28] ^ x[2];
  assign t[21] = t[29] ^ x[3];
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[6];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[9];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[29] = (x[1]);
  assign t[2] = ~(t[3] & t[9]);
  assign t[30] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[4]);
  assign t[32] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[7]);
  assign t[34] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[10]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[7] = ~(t[9] & t[8]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind21(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind22(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind23(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind24(x, y);
 input [12:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[3];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[9];
  assign t[15] = t[19] ^ x[12];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[8] ^ t[2];
  assign t[20] = t[28] ^ x[2];
  assign t[21] = t[29] ^ x[3];
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[6];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[9];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[29] = (x[1]);
  assign t[2] = ~(t[3] & t[9]);
  assign t[30] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[4]);
  assign t[32] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[7]);
  assign t[34] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[10]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[7] = ~(t[9] & t[8]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [12:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[3];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[21] & t[22]);
  assign t[17] = (~t[23] & t[24]);
  assign t[18] = (~t[25] & t[26]);
  assign t[19] = t[27] ^ x[2];
  assign t[1] = ~(t[7] ^ t[2]);
  assign t[20] = t[28] ^ x[3];
  assign t[21] = t[29] ^ x[5];
  assign t[22] = t[30] ^ x[6];
  assign t[23] = t[31] ^ x[8];
  assign t[24] = t[32] ^ x[9];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[12];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[1]);
  assign t[29] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[31] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[7]);
  assign t[33] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[10]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[6] = ~(t[7] & t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind28(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind29(x, y);
 input [12:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[3];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[21] & t[22]);
  assign t[17] = (~t[23] & t[24]);
  assign t[18] = (~t[25] & t[26]);
  assign t[19] = t[27] ^ x[2];
  assign t[1] = ~(t[7] ^ t[2]);
  assign t[20] = t[28] ^ x[3];
  assign t[21] = t[29] ^ x[5];
  assign t[22] = t[30] ^ x[6];
  assign t[23] = t[31] ^ x[8];
  assign t[24] = t[32] ^ x[9];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[12];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[1]);
  assign t[29] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[31] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[7]);
  assign t[33] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[10]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[6] = ~(t[7] & t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind31(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind32(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind33(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind34(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind36(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind37(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind38(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind39(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind41(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind46(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind51(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind56(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind61(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind66(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind71(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind76(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind81(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind86(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind91(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind96(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind101(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [16:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[11] ^ t[12];
  assign t[11] = x[11] ^ x[12];
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[28] & t[6]);
  assign t[14] = ~(t[30] & t[15]);
  assign t[15] = ~(t[29] & t[5]);
  assign t[16] = t[17] ^ t[18];
  assign t[17] = x[13] ^ x[14];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[6] & t[8]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = ~(t[21] & t[27]);
  assign t[21] = ~(t[22] & t[5]);
  assign t[22] = ~(t[30] & t[29]);
  assign t[23] = t[24] ^ t[25];
  assign t[24] = x[15] ^ x[16];
  assign t[25] = ~(t[19] & t[26]);
  assign t[26] = t[3] | t[27];
  assign t[27] = (t[31]);
  assign t[28] = (t[32]);
  assign t[29] = (t[33]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (t[34]);
  assign t[31] = t[35] ^ x[7];
  assign t[32] = t[36] ^ x[8];
  assign t[33] = t[37] ^ x[9];
  assign t[34] = t[38] ^ x[10];
  assign t[35] = (~t[39] & t[40]);
  assign t[36] = (~t[39] & t[41]);
  assign t[37] = (~t[39] & t[42]);
  assign t[38] = (~t[39] & t[43]);
  assign t[39] = t[44] ^ x[6];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[7];
  assign t[41] = t[46] ^ x[8];
  assign t[42] = t[47] ^ x[9];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[45] = (x[3]);
  assign t[46] = (x[4]);
  assign t[47] = (x[5]);
  assign t[48] = (x[2]);
  assign t[4] = ~(t[27] | t[7]);
  assign t[5] = ~(t[28]);
  assign t[6] = ~(t[29]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[30]);
  assign t[9] = ~(t[28] | t[29]);
  assign y = (t[0] & ~t[10] & ~t[16] & ~t[23]) | (~t[0] & t[10] & ~t[16] & ~t[23]) | (~t[0] & ~t[10] & t[16] & ~t[23]) | (~t[0] & ~t[10] & ~t[16] & t[23]) | (t[0] & t[10] & t[16] & ~t[23]) | (t[0] & t[10] & ~t[16] & t[23]) | (t[0] & ~t[10] & t[16] & t[23]) | (~t[0] & t[10] & t[16] & t[23]);
endmodule

module R2ind106(x, y);
 input [10:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[10];
  assign t[17] = (~t[21] & t[22]);
  assign t[18] = (~t[21] & t[23]);
  assign t[19] = (~t[21] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[21] & t[25]);
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = t[29] ^ x[9];
  assign t[25] = t[30] ^ x[10];
  assign t[26] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[27] = (x[3]);
  assign t[28] = (x[5]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = t[7] | t[9];
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[8] | t[5]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[2]);
  assign t[31] = (x[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[7] & t[10]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[12] & t[11]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [9:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[13]);
  assign t[11] = t[14] ^ x[7];
  assign t[12] = t[15] ^ x[8];
  assign t[13] = t[16] ^ x[9];
  assign t[14] = (~t[17] & t[18]);
  assign t[15] = (~t[17] & t[19]);
  assign t[16] = (~t[17] & t[20]);
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = t[23] ^ x[8];
  assign t[1] = x[0] ^ x[1];
  assign t[20] = t[24] ^ x[9];
  assign t[21] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[22] = (x[4]);
  assign t[23] = (x[2]);
  assign t[24] = (x[5]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[8] & t[5]);
  assign t[4] = ~(t[9] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[10] & t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = (t[11]);
  assign t[9] = (t[12]);
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [10:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[10];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[22] & t[24]);
  assign t[1] = x[0] ^ x[1];
  assign t[20] = (~t[22] & t[25]);
  assign t[21] = (~t[22] & t[26]);
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = t[30] ^ x[9];
  assign t[26] = t[31] ^ x[10];
  assign t[27] = (x[2] & ~x[3] & ~x[4] & ~x[5]) | (~x[2] & x[3] & ~x[4] & ~x[5]) | (~x[2] & ~x[3] & x[4] & ~x[5]) | (~x[2] & ~x[3] & ~x[4] & x[5]) | (x[2] & x[3] & x[4] & ~x[5]) | (x[2] & x[3] & ~x[4] & x[5]) | (x[2] & ~x[3] & x[4] & x[5]) | (~x[2] & x[3] & x[4] & x[5]);
  assign t[28] = (x[3]);
  assign t[29] = (x[4]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[5]);
  assign t[31] = (x[2]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(t[10] | t[7]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[13]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [163:0] x;
 output y;

 wire [635:0] t;
  assign t[0] = t[1] ? t[2] : t[388];
  assign t[100] = ~(t[410]);
  assign t[101] = ~(t[399] | t[400]);
  assign t[102] = ~(t[411]);
  assign t[103] = ~(t[412]);
  assign t[104] = ~(t[142] | t[143]);
  assign t[105] = ~(t[144] | t[145]);
  assign t[106] = ~(t[413]);
  assign t[107] = ~(t[414]);
  assign t[108] = ~(t[146] | t[147]);
  assign t[109] = ~(t[148] | t[149]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[415] | t[150]);
  assign t[111] = t[151] ? x[100] : x[99];
  assign t[112] = ~(t[152] & t[153]);
  assign t[113] = ~(t[416]);
  assign t[114] = ~(t[417]);
  assign t[115] = ~(t[154] | t[155]);
  assign t[116] = t[391] ? x[104] : x[103];
  assign t[117] = t[156] | t[157];
  assign t[118] = ~(t[391]);
  assign t[119] = ~(t[158] & t[392]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[159] & t[160]);
  assign t[121] = ~(t[77] | t[161]);
  assign t[122] = ~(t[77] | t[162]);
  assign t[123] = t[392] & t[163];
  assign t[124] = t[159] | t[158];
  assign t[125] = ~(t[164] & t[160]);
  assign t[126] = ~(x[7] & t[165]);
  assign t[127] = ~(t[159] & t[392]);
  assign t[128] = ~(t[158] & t[160]);
  assign t[129] = ~(t[391]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[140]);
  assign t[131] = ~(t[418]);
  assign t[132] = ~(t[405] | t[406]);
  assign t[133] = ~(t[166] | t[144]);
  assign t[134] = ~(t[167] | t[168]);
  assign t[135] = ~(t[419]);
  assign t[136] = ~(t[407] | t[408]);
  assign t[137] = ~(t[420]);
  assign t[138] = ~(t[421]);
  assign t[139] = ~(t[169] | t[170]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[171] | t[144]);
  assign t[141] = ~(t[172] | t[173]);
  assign t[142] = ~(t[422]);
  assign t[143] = ~(t[411] | t[412]);
  assign t[144] = ~(t[118] | t[174]);
  assign t[145] = t[175] | t[176];
  assign t[146] = ~(t[423]);
  assign t[147] = ~(t[413] | t[414]);
  assign t[148] = ~(t[424]);
  assign t[149] = ~(t[425]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[177] | t[178]);
  assign t[151] = ~(t[129]);
  assign t[152] = ~(t[156] | t[179]);
  assign t[153] = ~(t[47]);
  assign t[154] = ~(t[426]);
  assign t[155] = ~(t[416] | t[417]);
  assign t[156] = ~(t[180] & t[181]);
  assign t[157] = ~(t[182] & t[86]);
  assign t[158] = x[7] & t[390];
  assign t[159] = ~(x[7] | t[390]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[392]);
  assign t[161] = t[389] ? t[119] : t[120];
  assign t[162] = t[389] ? t[184] : t[183];
  assign t[163] = ~(t[118] | t[389]);
  assign t[164] = ~(x[7] | t[185]);
  assign t[165] = ~(t[390] | t[160]);
  assign t[166] = ~(t[118] | t[186]);
  assign t[167] = ~(t[31]);
  assign t[168] = ~(t[77] | t[187]);
  assign t[169] = ~(t[427]);
  assign t[16] = ~(t[389] & t[390]);
  assign t[170] = ~(t[420] | t[421]);
  assign t[171] = ~(t[118] | t[188]);
  assign t[172] = ~(t[189] & t[190]);
  assign t[173] = ~(t[80] & t[191]);
  assign t[174] = t[389] ? t[125] : t[184];
  assign t[175] = ~(t[77] | t[192]);
  assign t[176] = ~(t[180]);
  assign t[177] = ~(t[428]);
  assign t[178] = ~(t[424] | t[425]);
  assign t[179] = ~(t[193] & t[191]);
  assign t[17] = ~(t[391] & t[392]);
  assign t[180] = ~(t[163] & t[194]);
  assign t[181] = ~(t[165] & t[195]);
  assign t[182] = ~(t[47] | t[175]);
  assign t[183] = ~(t[392] & t[164]);
  assign t[184] = ~(x[7] & t[196]);
  assign t[185] = ~(t[390]);
  assign t[186] = t[389] ? t[120] : t[128];
  assign t[187] = t[389] ? t[183] : t[184];
  assign t[188] = t[389] ? t[128] : t[120];
  assign t[189] = ~(t[166] | t[197]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[118] & t[198]);
  assign t[191] = t[118] | t[199];
  assign t[192] = t[389] ? t[127] : t[128];
  assign t[193] = ~(t[144]);
  assign t[194] = ~(t[183] & t[126]);
  assign t[195] = t[77] & t[389];
  assign t[196] = ~(t[390] | t[392]);
  assign t[197] = ~(t[77] | t[200]);
  assign t[198] = ~(t[184] & t[183]);
  assign t[199] = t[389] ? t[184] : t[125];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[389] ? t[125] : t[126];
  assign t[201] = t[6] ? t[202] : t[429];
  assign t[202] = x[6] ? t[204] : t[203];
  assign t[203] = x[7] ? t[206] : t[205];
  assign t[204] = t[207] ^ x[117];
  assign t[205] = t[208] ^ t[209];
  assign t[206] = ~(t[210] ^ t[211]);
  assign t[207] = x[118] ^ x[119];
  assign t[208] = t[391] ? x[118] : x[119];
  assign t[209] = ~(t[212] ^ t[213]);
  assign t[20] = t[391] ? x[9] : x[10];
  assign t[210] = x[7] ? t[215] : t[214];
  assign t[211] = ~(t[216] ^ t[217]);
  assign t[212] = x[7] ? t[219] : t[218];
  assign t[213] = ~(t[220] ^ t[221]);
  assign t[214] = ~(t[222] & t[223]);
  assign t[215] = t[224] ^ t[218];
  assign t[216] = x[7] ? t[226] : t[225];
  assign t[217] = x[7] ? t[228] : t[227];
  assign t[218] = ~(t[229] & t[230]);
  assign t[219] = t[231] ^ t[232];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = x[7] ? t[234] : t[233];
  assign t[221] = x[7] ? t[236] : t[235];
  assign t[222] = ~(t[395] & t[52]);
  assign t[223] = ~(t[404] & t[237]);
  assign t[224] = t[85] ? x[121] : x[120];
  assign t[225] = ~(t[238] & t[239]);
  assign t[226] = t[240] ^ t[241];
  assign t[227] = ~(t[242] & t[243]);
  assign t[228] = t[244] ^ t[227];
  assign t[229] = ~(t[399] & t[64]);
  assign t[22] = ~(t[32] | t[33]);
  assign t[230] = ~(t[410] & t[245]);
  assign t[231] = t[85] ? x[123] : x[122];
  assign t[232] = ~(t[246] & t[247]);
  assign t[233] = ~(t[248] & t[249]);
  assign t[234] = t[250] ^ t[233];
  assign t[235] = ~(t[251] & t[252]);
  assign t[236] = t[253] ^ t[254];
  assign t[237] = ~(t[396] & t[51]);
  assign t[238] = ~(t[407] & t[94]);
  assign t[239] = ~(t[419] & t[255]);
  assign t[23] = ~(t[26] ^ t[34]);
  assign t[240] = t[85] ? x[125] : x[124];
  assign t[241] = ~(t[256] & t[257]);
  assign t[242] = ~(t[405] & t[89]);
  assign t[243] = ~(t[418] & t[258]);
  assign t[244] = t[85] ? x[127] : x[126];
  assign t[245] = ~(t[400] & t[63]);
  assign t[246] = ~(t[411] & t[103]);
  assign t[247] = ~(t[422] & t[259]);
  assign t[248] = ~(t[416] & t[114]);
  assign t[249] = ~(t[426] & t[260]);
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = t[391] ? x[129] : x[128];
  assign t[251] = ~(t[413] & t[107]);
  assign t[252] = ~(t[423] & t[261]);
  assign t[253] = t[391] ? x[131] : x[130];
  assign t[254] = ~(t[262] & t[263]);
  assign t[255] = ~(t[408] & t[93]);
  assign t[256] = ~(t[420] & t[138]);
  assign t[257] = ~(t[427] & t[264]);
  assign t[258] = ~(t[406] & t[88]);
  assign t[259] = ~(t[412] & t[102]);
  assign t[25] = x[7] ? t[38] : t[37];
  assign t[260] = ~(t[417] & t[113]);
  assign t[261] = ~(t[414] & t[106]);
  assign t[262] = ~(t[424] & t[149]);
  assign t[263] = ~(t[428] & t[265]);
  assign t[264] = ~(t[421] & t[137]);
  assign t[265] = ~(t[425] & t[148]);
  assign t[266] = t[1] ? t[267] : t[430];
  assign t[267] = x[6] ? t[269] : t[268];
  assign t[268] = x[7] ? t[271] : t[270];
  assign t[269] = t[272] ^ x[133];
  assign t[26] = ~(t[39] | t[40]);
  assign t[270] = t[273] ^ t[274];
  assign t[271] = ~(t[275] ^ t[276]);
  assign t[272] = x[134] ^ x[135];
  assign t[273] = t[391] ? x[134] : x[135];
  assign t[274] = ~(t[277] ^ t[278]);
  assign t[275] = x[7] ? t[280] : t[279];
  assign t[276] = ~(t[281] ^ t[282]);
  assign t[277] = x[7] ? t[284] : t[283];
  assign t[278] = ~(t[285] ^ t[286]);
  assign t[279] = ~(t[287] & t[288]);
  assign t[27] = ~(t[41] ^ t[42]);
  assign t[280] = t[289] ^ t[283];
  assign t[281] = x[7] ? t[291] : t[290];
  assign t[282] = x[7] ? t[293] : t[292];
  assign t[283] = ~(t[294] & t[295]);
  assign t[284] = t[296] ^ t[297];
  assign t[285] = x[7] ? t[299] : t[298];
  assign t[286] = x[7] ? t[301] : t[300];
  assign t[287] = ~(t[52] & t[83]);
  assign t[288] = ~(t[302] & t[393]);
  assign t[289] = t[85] ? x[137] : x[136];
  assign t[28] = x[7] ? t[44] : t[43];
  assign t[290] = ~(t[303] & t[304]);
  assign t[291] = t[305] ^ t[290];
  assign t[292] = ~(t[306] & t[307]);
  assign t[293] = t[308] ^ t[309];
  assign t[294] = ~(t[64] & t[100]);
  assign t[295] = ~(t[310] & t[394]);
  assign t[296] = t[311] ? x[139] : x[138];
  assign t[297] = ~(t[312] & t[313]);
  assign t[298] = ~(t[314] & t[315]);
  assign t[299] = t[316] ^ t[317];
  assign t[29] = x[7] ? t[46] : t[45];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = ~(t[318] & t[319]);
  assign t[301] = t[320] ^ t[300];
  assign t[302] = ~(t[321] & t[51]);
  assign t[303] = ~(t[89] & t[131]);
  assign t[304] = ~(t[322] & t[397]);
  assign t[305] = t[85] ? x[141] : x[140];
  assign t[306] = ~(t[94] & t[135]);
  assign t[307] = ~(t[323] & t[398]);
  assign t[308] = t[85] ? x[143] : x[142];
  assign t[309] = ~(t[324] & t[325]);
  assign t[30] = ~(t[47] | t[48]);
  assign t[310] = ~(t[326] & t[63]);
  assign t[311] = ~(t[129]);
  assign t[312] = ~(t[103] & t[142]);
  assign t[313] = ~(t[327] & t[401]);
  assign t[314] = ~(t[107] & t[146]);
  assign t[315] = ~(t[328] & t[402]);
  assign t[316] = t[391] ? x[145] : x[144];
  assign t[317] = ~(t[329] & t[330]);
  assign t[318] = ~(t[114] & t[154]);
  assign t[319] = ~(t[331] & t[403]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = t[391] ? x[147] : x[146];
  assign t[321] = ~(t[404] & t[396]);
  assign t[322] = ~(t[332] & t[88]);
  assign t[323] = ~(t[333] & t[93]);
  assign t[324] = ~(t[138] & t[169]);
  assign t[325] = ~(t[334] & t[409]);
  assign t[326] = ~(t[410] & t[400]);
  assign t[327] = ~(t[335] & t[102]);
  assign t[328] = ~(t[336] & t[106]);
  assign t[329] = ~(t[149] & t[177]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = ~(t[337] & t[415]);
  assign t[331] = ~(t[338] & t[113]);
  assign t[332] = ~(t[418] & t[406]);
  assign t[333] = ~(t[419] & t[408]);
  assign t[334] = ~(t[339] & t[137]);
  assign t[335] = ~(t[422] & t[412]);
  assign t[336] = ~(t[423] & t[414]);
  assign t[337] = ~(t[340] & t[148]);
  assign t[338] = ~(t[426] & t[417]);
  assign t[339] = ~(t[427] & t[421]);
  assign t[33] = ~(t[393] | t[53]);
  assign t[340] = ~(t[428] & t[425]);
  assign t[341] = t[6] ? t[342] : t[431];
  assign t[342] = x[6] ? t[344] : t[343];
  assign t[343] = x[7] ? t[346] : t[345];
  assign t[344] = t[347] ^ x[149];
  assign t[345] = t[348] ^ t[349];
  assign t[346] = ~(t[350] ^ t[351]);
  assign t[347] = x[150] ^ x[151];
  assign t[348] = t[391] ? x[150] : x[151];
  assign t[349] = ~(t[352] ^ t[353]);
  assign t[34] = ~(t[54] ^ t[55]);
  assign t[350] = x[7] ? t[355] : t[354];
  assign t[351] = ~(t[356] ^ t[357]);
  assign t[352] = x[7] ? t[359] : t[358];
  assign t[353] = ~(t[360] ^ t[361]);
  assign t[354] = ~(t[287] & t[362]);
  assign t[355] = t[363] ^ t[358];
  assign t[356] = x[7] ? t[365] : t[364];
  assign t[357] = x[7] ? t[367] : t[366];
  assign t[358] = ~(t[294] & t[368]);
  assign t[359] = t[369] ^ t[370];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = x[7] ? t[372] : t[371];
  assign t[361] = x[7] ? t[374] : t[373];
  assign t[362] = t[32] | t[393];
  assign t[363] = t[85] ? x[153] : x[152];
  assign t[364] = ~(t[303] & t[375]);
  assign t[365] = t[376] ^ t[364];
  assign t[366] = ~(t[306] & t[377]);
  assign t[367] = t[378] ^ t[379];
  assign t[368] = t[39] | t[394];
  assign t[369] = t[151] ? x[155] : x[154];
  assign t[36] = ~(t[35] ^ t[58]);
  assign t[370] = ~(t[312] & t[380]);
  assign t[371] = ~(t[314] & t[381]);
  assign t[372] = t[382] ^ t[383];
  assign t[373] = ~(t[318] & t[384]);
  assign t[374] = t[385] ^ t[373];
  assign t[375] = t[56] | t[397];
  assign t[376] = t[85] ? x[157] : x[156];
  assign t[377] = t[59] | t[398];
  assign t[378] = t[85] ? x[159] : x[158];
  assign t[379] = ~(t[324] & t[386]);
  assign t[37] = ~(t[59] | t[60]);
  assign t[380] = t[66] | t[401];
  assign t[381] = t[70] | t[402];
  assign t[382] = t[391] ? x[161] : x[160];
  assign t[383] = ~(t[329] & t[387]);
  assign t[384] = t[74] | t[403];
  assign t[385] = t[391] ? x[163] : x[162];
  assign t[386] = t[96] | t[409];
  assign t[387] = t[109] | t[415];
  assign t[388] = (t[432]);
  assign t[389] = (t[433]);
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = (t[434]);
  assign t[391] = (t[435]);
  assign t[392] = (t[436]);
  assign t[393] = (t[437]);
  assign t[394] = (t[438]);
  assign t[395] = (t[439]);
  assign t[396] = (t[440]);
  assign t[397] = (t[441]);
  assign t[398] = (t[442]);
  assign t[399] = (t[443]);
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (t[444]);
  assign t[401] = (t[445]);
  assign t[402] = (t[446]);
  assign t[403] = (t[447]);
  assign t[404] = (t[448]);
  assign t[405] = (t[449]);
  assign t[406] = (t[450]);
  assign t[407] = (t[451]);
  assign t[408] = (t[452]);
  assign t[409] = (t[453]);
  assign t[40] = ~(t[394] | t[65]);
  assign t[410] = (t[454]);
  assign t[411] = (t[455]);
  assign t[412] = (t[456]);
  assign t[413] = (t[457]);
  assign t[414] = (t[458]);
  assign t[415] = (t[459]);
  assign t[416] = (t[460]);
  assign t[417] = (t[461]);
  assign t[418] = (t[462]);
  assign t[419] = (t[463]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (t[464]);
  assign t[421] = (t[465]);
  assign t[422] = (t[466]);
  assign t[423] = (t[467]);
  assign t[424] = (t[468]);
  assign t[425] = (t[469]);
  assign t[426] = (t[470]);
  assign t[427] = (t[471]);
  assign t[428] = (t[472]);
  assign t[429] = (t[473]);
  assign t[42] = ~(t[68] ^ t[69]);
  assign t[430] = (t[474]);
  assign t[431] = (t[475]);
  assign t[432] = t[476] ^ x[5];
  assign t[433] = t[477] ^ x[13];
  assign t[434] = t[478] ^ x[16];
  assign t[435] = t[479] ^ x[19];
  assign t[436] = t[480] ^ x[22];
  assign t[437] = t[481] ^ x[28];
  assign t[438] = t[482] ^ x[34];
  assign t[439] = t[483] ^ x[35];
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = t[484] ^ x[36];
  assign t[441] = t[485] ^ x[44];
  assign t[442] = t[486] ^ x[50];
  assign t[443] = t[487] ^ x[51];
  assign t[444] = t[488] ^ x[52];
  assign t[445] = t[489] ^ x[58];
  assign t[446] = t[490] ^ x[66];
  assign t[447] = t[491] ^ x[72];
  assign t[448] = t[492] ^ x[73];
  assign t[449] = t[493] ^ x[74];
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = t[494] ^ x[75];
  assign t[451] = t[495] ^ x[78];
  assign t[452] = t[496] ^ x[79];
  assign t[453] = t[497] ^ x[85];
  assign t[454] = t[498] ^ x[88];
  assign t[455] = t[499] ^ x[89];
  assign t[456] = t[500] ^ x[90];
  assign t[457] = t[501] ^ x[91];
  assign t[458] = t[502] ^ x[92];
  assign t[459] = t[503] ^ x[98];
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = t[504] ^ x[101];
  assign t[461] = t[505] ^ x[102];
  assign t[462] = t[506] ^ x[105];
  assign t[463] = t[507] ^ x[106];
  assign t[464] = t[508] ^ x[107];
  assign t[465] = t[509] ^ x[108];
  assign t[466] = t[510] ^ x[109];
  assign t[467] = t[511] ^ x[110];
  assign t[468] = t[512] ^ x[111];
  assign t[469] = t[513] ^ x[112];
  assign t[46] = ~(t[45] ^ t[76]);
  assign t[470] = t[514] ^ x[113];
  assign t[471] = t[515] ^ x[114];
  assign t[472] = t[516] ^ x[115];
  assign t[473] = t[517] ^ x[116];
  assign t[474] = t[518] ^ x[132];
  assign t[475] = t[519] ^ x[148];
  assign t[476] = (~t[520] & t[521]);
  assign t[477] = (~t[522] & t[523]);
  assign t[478] = (~t[524] & t[525]);
  assign t[479] = (~t[526] & t[527]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = (~t[528] & t[529]);
  assign t[481] = (~t[530] & t[531]);
  assign t[482] = (~t[532] & t[533]);
  assign t[483] = (~t[530] & t[534]);
  assign t[484] = (~t[530] & t[535]);
  assign t[485] = (~t[536] & t[537]);
  assign t[486] = (~t[538] & t[539]);
  assign t[487] = (~t[532] & t[540]);
  assign t[488] = (~t[532] & t[541]);
  assign t[489] = (~t[542] & t[543]);
  assign t[48] = ~(t[79] & t[80]);
  assign t[490] = (~t[544] & t[545]);
  assign t[491] = (~t[546] & t[547]);
  assign t[492] = (~t[530] & t[548]);
  assign t[493] = (~t[536] & t[549]);
  assign t[494] = (~t[536] & t[550]);
  assign t[495] = (~t[538] & t[551]);
  assign t[496] = (~t[538] & t[552]);
  assign t[497] = (~t[553] & t[554]);
  assign t[498] = (~t[532] & t[555]);
  assign t[499] = (~t[542] & t[556]);
  assign t[49] = ~(t[77] | t[81]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[542] & t[557]);
  assign t[501] = (~t[544] & t[558]);
  assign t[502] = (~t[544] & t[559]);
  assign t[503] = (~t[560] & t[561]);
  assign t[504] = (~t[546] & t[562]);
  assign t[505] = (~t[546] & t[563]);
  assign t[506] = (~t[536] & t[564]);
  assign t[507] = (~t[538] & t[565]);
  assign t[508] = (~t[553] & t[566]);
  assign t[509] = (~t[553] & t[567]);
  assign t[50] = ~(t[77] | t[82]);
  assign t[510] = (~t[542] & t[568]);
  assign t[511] = (~t[544] & t[569]);
  assign t[512] = (~t[560] & t[570]);
  assign t[513] = (~t[560] & t[571]);
  assign t[514] = (~t[546] & t[572]);
  assign t[515] = (~t[553] & t[573]);
  assign t[516] = (~t[560] & t[574]);
  assign t[517] = (~t[520] & t[575]);
  assign t[518] = (~t[520] & t[576]);
  assign t[519] = (~t[520] & t[577]);
  assign t[51] = ~(t[395]);
  assign t[520] = t[578] ^ x[4];
  assign t[521] = t[579] ^ x[5];
  assign t[522] = t[580] ^ x[12];
  assign t[523] = t[581] ^ x[13];
  assign t[524] = t[582] ^ x[15];
  assign t[525] = t[583] ^ x[16];
  assign t[526] = t[584] ^ x[18];
  assign t[527] = t[585] ^ x[19];
  assign t[528] = t[586] ^ x[21];
  assign t[529] = t[587] ^ x[22];
  assign t[52] = ~(t[396]);
  assign t[530] = t[588] ^ x[27];
  assign t[531] = t[589] ^ x[28];
  assign t[532] = t[590] ^ x[33];
  assign t[533] = t[591] ^ x[34];
  assign t[534] = t[592] ^ x[35];
  assign t[535] = t[593] ^ x[36];
  assign t[536] = t[594] ^ x[43];
  assign t[537] = t[595] ^ x[44];
  assign t[538] = t[596] ^ x[49];
  assign t[539] = t[597] ^ x[50];
  assign t[53] = ~(t[83] | t[84]);
  assign t[540] = t[598] ^ x[51];
  assign t[541] = t[599] ^ x[52];
  assign t[542] = t[600] ^ x[57];
  assign t[543] = t[601] ^ x[58];
  assign t[544] = t[602] ^ x[65];
  assign t[545] = t[603] ^ x[66];
  assign t[546] = t[604] ^ x[71];
  assign t[547] = t[605] ^ x[72];
  assign t[548] = t[606] ^ x[73];
  assign t[549] = t[607] ^ x[74];
  assign t[54] = t[85] ? x[38] : x[37];
  assign t[550] = t[608] ^ x[75];
  assign t[551] = t[609] ^ x[78];
  assign t[552] = t[610] ^ x[79];
  assign t[553] = t[611] ^ x[84];
  assign t[554] = t[612] ^ x[85];
  assign t[555] = t[613] ^ x[88];
  assign t[556] = t[614] ^ x[89];
  assign t[557] = t[615] ^ x[90];
  assign t[558] = t[616] ^ x[91];
  assign t[559] = t[617] ^ x[92];
  assign t[55] = ~(t[86] & t[87]);
  assign t[560] = t[618] ^ x[97];
  assign t[561] = t[619] ^ x[98];
  assign t[562] = t[620] ^ x[101];
  assign t[563] = t[621] ^ x[102];
  assign t[564] = t[622] ^ x[105];
  assign t[565] = t[623] ^ x[106];
  assign t[566] = t[624] ^ x[107];
  assign t[567] = t[625] ^ x[108];
  assign t[568] = t[626] ^ x[109];
  assign t[569] = t[627] ^ x[110];
  assign t[56] = ~(t[88] | t[89]);
  assign t[570] = t[628] ^ x[111];
  assign t[571] = t[629] ^ x[112];
  assign t[572] = t[630] ^ x[113];
  assign t[573] = t[631] ^ x[114];
  assign t[574] = t[632] ^ x[115];
  assign t[575] = t[633] ^ x[116];
  assign t[576] = t[634] ^ x[132];
  assign t[577] = t[635] ^ x[148];
  assign t[578] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[579] = (x[0]);
  assign t[57] = ~(t[397] | t[90]);
  assign t[580] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[581] = (x[11]);
  assign t[582] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[583] = (x[14]);
  assign t[584] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[585] = (x[17]);
  assign t[586] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[587] = (x[20]);
  assign t[588] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[589] = (x[24]);
  assign t[58] = ~(t[91] ^ t[92]);
  assign t[590] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[591] = (x[30]);
  assign t[592] = (x[25]);
  assign t[593] = (x[26]);
  assign t[594] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[595] = (x[40]);
  assign t[596] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[597] = (x[46]);
  assign t[598] = (x[31]);
  assign t[599] = (x[32]);
  assign t[59] = ~(t[93] | t[94]);
  assign t[5] = t[9] ^ x[8];
  assign t[600] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[601] = (x[54]);
  assign t[602] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[603] = (x[62]);
  assign t[604] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[605] = (x[68]);
  assign t[606] = (x[23]);
  assign t[607] = (x[41]);
  assign t[608] = (x[42]);
  assign t[609] = (x[47]);
  assign t[60] = ~(t[398] | t[95]);
  assign t[610] = (x[48]);
  assign t[611] = (x[80] & ~x[81] & ~x[82] & ~x[83]) | (~x[80] & x[81] & ~x[82] & ~x[83]) | (~x[80] & ~x[81] & x[82] & ~x[83]) | (~x[80] & ~x[81] & ~x[82] & x[83]) | (x[80] & x[81] & x[82] & ~x[83]) | (x[80] & x[81] & ~x[82] & x[83]) | (x[80] & ~x[81] & x[82] & x[83]) | (~x[80] & x[81] & x[82] & x[83]);
  assign t[612] = (x[81]);
  assign t[613] = (x[29]);
  assign t[614] = (x[55]);
  assign t[615] = (x[56]);
  assign t[616] = (x[63]);
  assign t[617] = (x[64]);
  assign t[618] = (x[93] & ~x[94] & ~x[95] & ~x[96]) | (~x[93] & x[94] & ~x[95] & ~x[96]) | (~x[93] & ~x[94] & x[95] & ~x[96]) | (~x[93] & ~x[94] & ~x[95] & x[96]) | (x[93] & x[94] & x[95] & ~x[96]) | (x[93] & x[94] & ~x[95] & x[96]) | (x[93] & ~x[94] & x[95] & x[96]) | (~x[93] & x[94] & x[95] & x[96]);
  assign t[619] = (x[94]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[620] = (x[69]);
  assign t[621] = (x[70]);
  assign t[622] = (x[39]);
  assign t[623] = (x[45]);
  assign t[624] = (x[82]);
  assign t[625] = (x[83]);
  assign t[626] = (x[53]);
  assign t[627] = (x[61]);
  assign t[628] = (x[95]);
  assign t[629] = (x[96]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[630] = (x[67]);
  assign t[631] = (x[80]);
  assign t[632] = (x[93]);
  assign t[633] = (x[1]);
  assign t[634] = (x[2]);
  assign t[635] = (x[3]);
  assign t[63] = ~(t[399]);
  assign t[64] = ~(t[400]);
  assign t[65] = ~(t[100] | t[101]);
  assign t[66] = ~(t[102] | t[103]);
  assign t[67] = ~(t[401] | t[104]);
  assign t[68] = t[391] ? x[60] : x[59];
  assign t[69] = ~(t[30] & t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[402] | t[108]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[111] ^ t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[403] | t[115]);
  assign t[76] = ~(t[116] ^ t[117]);
  assign t[77] = ~(t[118]);
  assign t[78] = t[389] ? t[120] : t[119];
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[123] & t[124]);
  assign t[81] = t[389] ? t[126] : t[125];
  assign t[82] = t[389] ? t[128] : t[127];
  assign t[83] = ~(t[404]);
  assign t[84] = ~(t[395] | t[396]);
  assign t[85] = ~(t[129]);
  assign t[86] = ~(t[122] | t[50]);
  assign t[87] = ~(t[123] | t[130]);
  assign t[88] = ~(t[405]);
  assign t[89] = ~(t[406]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = t[85] ? x[77] : x[76];
  assign t[92] = ~(t[133] & t[134]);
  assign t[93] = ~(t[407]);
  assign t[94] = ~(t[408]);
  assign t[95] = ~(t[135] | t[136]);
  assign t[96] = ~(t[137] | t[138]);
  assign t[97] = ~(t[409] | t[139]);
  assign t[98] = t[85] ? x[87] : x[86];
  assign t[99] = ~(t[140] & t[141]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[201] & ~t[266] & ~t[341]) | (~t[0] & t[201] & ~t[266] & ~t[341]) | (~t[0] & ~t[201] & t[266] & ~t[341]) | (~t[0] & ~t[201] & ~t[266] & t[341]) | (t[0] & t[201] & t[266] & ~t[341]) | (t[0] & t[201] & ~t[266] & t[341]) | (t[0] & ~t[201] & t[266] & t[341]) | (~t[0] & t[201] & t[266] & t[341]);
endmodule

module R2ind111(x, y);
 input [115:0] x;
 output y;

 wire [332:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[141]);
  assign t[101] = (t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[103] ? x[21] : x[22];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = t[182] ^ x[5];
  assign t[142] = t[183] ^ x[11];
  assign t[143] = t[184] ^ x[14];
  assign t[144] = t[185] ^ x[17];
  assign t[145] = t[186] ^ x[20];
  assign t[146] = t[187] ^ x[28];
  assign t[147] = t[188] ^ x[36];
  assign t[148] = t[189] ^ x[39];
  assign t[149] = t[190] ^ x[40];
  assign t[14] = x[7] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[46];
  assign t[151] = t[192] ^ x[54];
  assign t[152] = t[193] ^ x[57];
  assign t[153] = t[194] ^ x[58];
  assign t[154] = t[195] ^ x[64];
  assign t[155] = t[196] ^ x[70];
  assign t[156] = t[197] ^ x[78];
  assign t[157] = t[198] ^ x[81];
  assign t[158] = t[199] ^ x[82];
  assign t[159] = t[200] ^ x[83];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[84];
  assign t[161] = t[202] ^ x[85];
  assign t[162] = t[203] ^ x[91];
  assign t[163] = t[204] ^ x[92];
  assign t[164] = t[205] ^ x[93];
  assign t[165] = t[206] ^ x[94];
  assign t[166] = t[207] ^ x[95];
  assign t[167] = t[208] ^ x[96];
  assign t[168] = t[209] ^ x[102];
  assign t[169] = t[210] ^ x[103];
  assign t[16] = x[7] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[104];
  assign t[171] = t[212] ^ x[105];
  assign t[172] = t[213] ^ x[106];
  assign t[173] = t[214] ^ x[107];
  assign t[174] = t[215] ^ x[108];
  assign t[175] = t[216] ^ x[109];
  assign t[176] = t[217] ^ x[110];
  assign t[177] = t[218] ^ x[111];
  assign t[178] = t[219] ^ x[112];
  assign t[179] = t[220] ^ x[113];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[114];
  assign t[181] = t[222] ^ x[115];
  assign t[182] = (~t[223] & t[224]);
  assign t[183] = (~t[225] & t[226]);
  assign t[184] = (~t[227] & t[228]);
  assign t[185] = (~t[229] & t[230]);
  assign t[186] = (~t[231] & t[232]);
  assign t[187] = (~t[233] & t[234]);
  assign t[188] = (~t[235] & t[236]);
  assign t[189] = (~t[233] & t[237]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (~t[233] & t[238]);
  assign t[191] = (~t[239] & t[240]);
  assign t[192] = (~t[241] & t[242]);
  assign t[193] = (~t[235] & t[243]);
  assign t[194] = (~t[235] & t[244]);
  assign t[195] = (~t[245] & t[246]);
  assign t[196] = (~t[247] & t[248]);
  assign t[197] = (~t[249] & t[250]);
  assign t[198] = (~t[233] & t[251]);
  assign t[199] = (~t[239] & t[252]);
  assign t[19] = t[28] ^ t[22];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (~t[239] & t[253]);
  assign t[201] = (~t[241] & t[254]);
  assign t[202] = (~t[241] & t[255]);
  assign t[203] = (~t[256] & t[257]);
  assign t[204] = (~t[235] & t[258]);
  assign t[205] = (~t[245] & t[259]);
  assign t[206] = (~t[245] & t[260]);
  assign t[207] = (~t[247] & t[261]);
  assign t[208] = (~t[247] & t[262]);
  assign t[209] = (~t[263] & t[264]);
  assign t[20] = x[7] ? t[30] : t[29];
  assign t[210] = (~t[249] & t[265]);
  assign t[211] = (~t[249] & t[266]);
  assign t[212] = (~t[239] & t[267]);
  assign t[213] = (~t[241] & t[268]);
  assign t[214] = (~t[256] & t[269]);
  assign t[215] = (~t[256] & t[270]);
  assign t[216] = (~t[245] & t[271]);
  assign t[217] = (~t[247] & t[272]);
  assign t[218] = (~t[263] & t[273]);
  assign t[219] = (~t[263] & t[274]);
  assign t[21] = x[7] ? t[32] : t[31];
  assign t[220] = (~t[249] & t[275]);
  assign t[221] = (~t[256] & t[276]);
  assign t[222] = (~t[263] & t[277]);
  assign t[223] = t[278] ^ x[4];
  assign t[224] = t[279] ^ x[5];
  assign t[225] = t[280] ^ x[10];
  assign t[226] = t[281] ^ x[11];
  assign t[227] = t[282] ^ x[13];
  assign t[228] = t[283] ^ x[14];
  assign t[229] = t[284] ^ x[16];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[285] ^ x[17];
  assign t[231] = t[286] ^ x[19];
  assign t[232] = t[287] ^ x[20];
  assign t[233] = t[288] ^ x[27];
  assign t[234] = t[289] ^ x[28];
  assign t[235] = t[290] ^ x[35];
  assign t[236] = t[291] ^ x[36];
  assign t[237] = t[292] ^ x[39];
  assign t[238] = t[293] ^ x[40];
  assign t[239] = t[294] ^ x[45];
  assign t[23] = t[35] ^ t[36];
  assign t[240] = t[295] ^ x[46];
  assign t[241] = t[296] ^ x[53];
  assign t[242] = t[297] ^ x[54];
  assign t[243] = t[298] ^ x[57];
  assign t[244] = t[299] ^ x[58];
  assign t[245] = t[300] ^ x[63];
  assign t[246] = t[301] ^ x[64];
  assign t[247] = t[302] ^ x[69];
  assign t[248] = t[303] ^ x[70];
  assign t[249] = t[304] ^ x[77];
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = t[305] ^ x[78];
  assign t[251] = t[306] ^ x[81];
  assign t[252] = t[307] ^ x[82];
  assign t[253] = t[308] ^ x[83];
  assign t[254] = t[309] ^ x[84];
  assign t[255] = t[310] ^ x[85];
  assign t[256] = t[311] ^ x[90];
  assign t[257] = t[312] ^ x[91];
  assign t[258] = t[313] ^ x[92];
  assign t[259] = t[314] ^ x[93];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[315] ^ x[94];
  assign t[261] = t[316] ^ x[95];
  assign t[262] = t[317] ^ x[96];
  assign t[263] = t[318] ^ x[101];
  assign t[264] = t[319] ^ x[102];
  assign t[265] = t[320] ^ x[103];
  assign t[266] = t[321] ^ x[104];
  assign t[267] = t[322] ^ x[105];
  assign t[268] = t[323] ^ x[106];
  assign t[269] = t[324] ^ x[107];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[325] ^ x[108];
  assign t[271] = t[326] ^ x[109];
  assign t[272] = t[327] ^ x[110];
  assign t[273] = t[328] ^ x[111];
  assign t[274] = t[329] ^ x[112];
  assign t[275] = t[330] ^ x[113];
  assign t[276] = t[331] ^ x[114];
  assign t[277] = t[332] ^ x[115];
  assign t[278] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[279] = (x[3]);
  assign t[27] = t[43] | t[105];
  assign t[280] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[281] = (x[9]);
  assign t[282] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[283] = (x[12]);
  assign t[284] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[285] = (x[15]);
  assign t[286] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[287] = (x[18]);
  assign t[288] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[289] = (x[24]);
  assign t[28] = t[44] ? x[30] : x[29];
  assign t[290] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[291] = (x[32]);
  assign t[292] = (x[26]);
  assign t[293] = (x[23]);
  assign t[294] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[295] = (x[42]);
  assign t[296] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[297] = (x[50]);
  assign t[298] = (x[34]);
  assign t[299] = (x[31]);
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[301] = (x[60]);
  assign t[302] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[303] = (x[66]);
  assign t[304] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[305] = (x[74]);
  assign t[306] = (x[25]);
  assign t[307] = (x[44]);
  assign t[308] = (x[41]);
  assign t[309] = (x[52]);
  assign t[30] = t[47] ^ t[29];
  assign t[310] = (x[49]);
  assign t[311] = (x[86] & ~x[87] & ~x[88] & ~x[89]) | (~x[86] & x[87] & ~x[88] & ~x[89]) | (~x[86] & ~x[87] & x[88] & ~x[89]) | (~x[86] & ~x[87] & ~x[88] & x[89]) | (x[86] & x[87] & x[88] & ~x[89]) | (x[86] & x[87] & ~x[88] & x[89]) | (x[86] & ~x[87] & x[88] & x[89]) | (~x[86] & x[87] & x[88] & x[89]);
  assign t[312] = (x[87]);
  assign t[313] = (x[33]);
  assign t[314] = (x[62]);
  assign t[315] = (x[59]);
  assign t[316] = (x[68]);
  assign t[317] = (x[65]);
  assign t[318] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[319] = (x[98]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = (x[76]);
  assign t[321] = (x[73]);
  assign t[322] = (x[43]);
  assign t[323] = (x[51]);
  assign t[324] = (x[89]);
  assign t[325] = (x[86]);
  assign t[326] = (x[61]);
  assign t[327] = (x[67]);
  assign t[328] = (x[100]);
  assign t[329] = (x[97]);
  assign t[32] = t[50] ^ t[51];
  assign t[330] = (x[75]);
  assign t[331] = (x[88]);
  assign t[332] = (x[99]);
  assign t[33] = ~(t[52] & t[53]);
  assign t[34] = t[54] | t[106];
  assign t[35] = t[55] ? x[38] : x[37];
  assign t[36] = ~(t[56] & t[57]);
  assign t[37] = ~(t[58] & t[59]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = ~(t[62] & t[63]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[64] ^ t[39];
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[108]);
  assign t[43] = ~(t[65] | t[41]);
  assign t[44] = ~(t[66]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = t[69] | t[109];
  assign t[47] = t[44] ? x[48] : x[47];
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = t[72] | t[110];
  assign t[4] = ~(x[6]);
  assign t[50] = t[44] ? x[56] : x[55];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[111]);
  assign t[53] = ~(t[112]);
  assign t[54] = ~(t[75] | t[52]);
  assign t[55] = ~(t[66]);
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = t[78] | t[113];
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = t[81] | t[114];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[103] ? x[72] : x[71];
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[115];
  assign t[64] = t[103] ? x[80] : x[79];
  assign t[65] = ~(t[116]);
  assign t[66] = ~(t[103]);
  assign t[67] = ~(t[117]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[87] | t[67]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[119]);
  assign t[71] = ~(t[120]);
  assign t[72] = ~(t[88] | t[70]);
  assign t[73] = ~(t[89] & t[90]);
  assign t[74] = t[91] | t[121];
  assign t[75] = ~(t[122]);
  assign t[76] = ~(t[123]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[92] | t[76]);
  assign t[79] = ~(t[125]);
  assign t[7] = ~(t[101] & t[102]);
  assign t[80] = ~(t[126]);
  assign t[81] = ~(t[93] | t[79]);
  assign t[82] = ~(t[94] & t[95]);
  assign t[83] = t[96] | t[127];
  assign t[84] = ~(t[128]);
  assign t[85] = ~(t[129]);
  assign t[86] = ~(t[97] | t[84]);
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[103] & t[104]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[98] | t[89]);
  assign t[92] = ~(t[134]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[99] | t[94]);
  assign t[97] = ~(t[138]);
  assign t[98] = ~(t[139]);
  assign t[99] = ~(t[140]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [115:0] x;
 output y;

 wire [343:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[109] & t[110]);
  assign t[105] = ~(t[140] & t[139]);
  assign t[106] = ~(t[149]);
  assign t[107] = ~(t[144] & t[143]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[148] & t[147]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[112] ? x[9] : x[10];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[7] ? t[21] : t[20];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[5];
  assign t[153] = t[194] ^ x[13];
  assign t[154] = t[195] ^ x[16];
  assign t[155] = t[196] ^ x[19];
  assign t[156] = t[197] ^ x[22];
  assign t[157] = t[198] ^ x[28];
  assign t[158] = t[199] ^ x[36];
  assign t[159] = t[200] ^ x[39];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[201] ^ x[40];
  assign t[161] = t[202] ^ x[46];
  assign t[162] = t[203] ^ x[54];
  assign t[163] = t[204] ^ x[57];
  assign t[164] = t[205] ^ x[58];
  assign t[165] = t[206] ^ x[64];
  assign t[166] = t[207] ^ x[70];
  assign t[167] = t[208] ^ x[78];
  assign t[168] = t[209] ^ x[81];
  assign t[169] = t[210] ^ x[82];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[83];
  assign t[171] = t[212] ^ x[84];
  assign t[172] = t[213] ^ x[85];
  assign t[173] = t[214] ^ x[91];
  assign t[174] = t[215] ^ x[92];
  assign t[175] = t[216] ^ x[93];
  assign t[176] = t[217] ^ x[94];
  assign t[177] = t[218] ^ x[95];
  assign t[178] = t[219] ^ x[96];
  assign t[179] = t[220] ^ x[102];
  assign t[17] = ~(t[112] & t[115]);
  assign t[180] = t[221] ^ x[103];
  assign t[181] = t[222] ^ x[104];
  assign t[182] = t[223] ^ x[105];
  assign t[183] = t[224] ^ x[106];
  assign t[184] = t[225] ^ x[107];
  assign t[185] = t[226] ^ x[108];
  assign t[186] = t[227] ^ x[109];
  assign t[187] = t[228] ^ x[110];
  assign t[188] = t[229] ^ x[111];
  assign t[189] = t[230] ^ x[112];
  assign t[18] = x[7] ? t[25] : t[24];
  assign t[190] = t[231] ^ x[113];
  assign t[191] = t[232] ^ x[114];
  assign t[192] = t[233] ^ x[115];
  assign t[193] = (~t[234] & t[235]);
  assign t[194] = (~t[236] & t[237]);
  assign t[195] = (~t[238] & t[239]);
  assign t[196] = (~t[240] & t[241]);
  assign t[197] = (~t[242] & t[243]);
  assign t[198] = (~t[244] & t[245]);
  assign t[199] = (~t[246] & t[247]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[244] & t[248]);
  assign t[201] = (~t[244] & t[249]);
  assign t[202] = (~t[250] & t[251]);
  assign t[203] = (~t[252] & t[253]);
  assign t[204] = (~t[246] & t[254]);
  assign t[205] = (~t[246] & t[255]);
  assign t[206] = (~t[256] & t[257]);
  assign t[207] = (~t[258] & t[259]);
  assign t[208] = (~t[260] & t[261]);
  assign t[209] = (~t[244] & t[262]);
  assign t[20] = ~(t[28] & t[29]);
  assign t[210] = (~t[250] & t[263]);
  assign t[211] = (~t[250] & t[264]);
  assign t[212] = (~t[252] & t[265]);
  assign t[213] = (~t[252] & t[266]);
  assign t[214] = (~t[267] & t[268]);
  assign t[215] = (~t[246] & t[269]);
  assign t[216] = (~t[256] & t[270]);
  assign t[217] = (~t[256] & t[271]);
  assign t[218] = (~t[258] & t[272]);
  assign t[219] = (~t[258] & t[273]);
  assign t[21] = t[30] ^ t[24];
  assign t[220] = (~t[274] & t[275]);
  assign t[221] = (~t[260] & t[276]);
  assign t[222] = (~t[260] & t[277]);
  assign t[223] = (~t[250] & t[278]);
  assign t[224] = (~t[252] & t[279]);
  assign t[225] = (~t[267] & t[280]);
  assign t[226] = (~t[267] & t[281]);
  assign t[227] = (~t[256] & t[282]);
  assign t[228] = (~t[258] & t[283]);
  assign t[229] = (~t[274] & t[284]);
  assign t[22] = x[7] ? t[32] : t[31];
  assign t[230] = (~t[274] & t[285]);
  assign t[231] = (~t[260] & t[286]);
  assign t[232] = (~t[267] & t[287]);
  assign t[233] = (~t[274] & t[288]);
  assign t[234] = t[289] ^ x[4];
  assign t[235] = t[290] ^ x[5];
  assign t[236] = t[291] ^ x[12];
  assign t[237] = t[292] ^ x[13];
  assign t[238] = t[293] ^ x[15];
  assign t[239] = t[294] ^ x[16];
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = t[295] ^ x[18];
  assign t[241] = t[296] ^ x[19];
  assign t[242] = t[297] ^ x[21];
  assign t[243] = t[298] ^ x[22];
  assign t[244] = t[299] ^ x[27];
  assign t[245] = t[300] ^ x[28];
  assign t[246] = t[301] ^ x[35];
  assign t[247] = t[302] ^ x[36];
  assign t[248] = t[303] ^ x[39];
  assign t[249] = t[304] ^ x[40];
  assign t[24] = ~(t[35] & t[36]);
  assign t[250] = t[305] ^ x[45];
  assign t[251] = t[306] ^ x[46];
  assign t[252] = t[307] ^ x[53];
  assign t[253] = t[308] ^ x[54];
  assign t[254] = t[309] ^ x[57];
  assign t[255] = t[310] ^ x[58];
  assign t[256] = t[311] ^ x[63];
  assign t[257] = t[312] ^ x[64];
  assign t[258] = t[313] ^ x[69];
  assign t[259] = t[314] ^ x[70];
  assign t[25] = t[37] ^ t[38];
  assign t[260] = t[315] ^ x[77];
  assign t[261] = t[316] ^ x[78];
  assign t[262] = t[317] ^ x[81];
  assign t[263] = t[318] ^ x[82];
  assign t[264] = t[319] ^ x[83];
  assign t[265] = t[320] ^ x[84];
  assign t[266] = t[321] ^ x[85];
  assign t[267] = t[322] ^ x[90];
  assign t[268] = t[323] ^ x[91];
  assign t[269] = t[324] ^ x[92];
  assign t[26] = x[7] ? t[40] : t[39];
  assign t[270] = t[325] ^ x[93];
  assign t[271] = t[326] ^ x[94];
  assign t[272] = t[327] ^ x[95];
  assign t[273] = t[328] ^ x[96];
  assign t[274] = t[329] ^ x[101];
  assign t[275] = t[330] ^ x[102];
  assign t[276] = t[331] ^ x[103];
  assign t[277] = t[332] ^ x[104];
  assign t[278] = t[333] ^ x[105];
  assign t[279] = t[334] ^ x[106];
  assign t[27] = x[7] ? t[42] : t[41];
  assign t[280] = t[335] ^ x[107];
  assign t[281] = t[336] ^ x[108];
  assign t[282] = t[337] ^ x[109];
  assign t[283] = t[338] ^ x[110];
  assign t[284] = t[339] ^ x[111];
  assign t[285] = t[340] ^ x[112];
  assign t[286] = t[341] ^ x[113];
  assign t[287] = t[342] ^ x[114];
  assign t[288] = t[343] ^ x[115];
  assign t[289] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = ~(t[43] & t[44]);
  assign t[290] = (x[2]);
  assign t[291] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[292] = (x[11]);
  assign t[293] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[294] = (x[14]);
  assign t[295] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[296] = (x[17]);
  assign t[297] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[298] = (x[20]);
  assign t[299] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[29] = ~(t[45] & t[116]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[24]);
  assign t[301] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[302] = (x[32]);
  assign t[303] = (x[26]);
  assign t[304] = (x[23]);
  assign t[305] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[306] = (x[42]);
  assign t[307] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[308] = (x[50]);
  assign t[309] = (x[34]);
  assign t[30] = t[46] ? x[30] : x[29];
  assign t[310] = (x[31]);
  assign t[311] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[312] = (x[60]);
  assign t[313] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[314] = (x[66]);
  assign t[315] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[316] = (x[74]);
  assign t[317] = (x[25]);
  assign t[318] = (x[44]);
  assign t[319] = (x[41]);
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = (x[52]);
  assign t[321] = (x[49]);
  assign t[322] = (x[86] & ~x[87] & ~x[88] & ~x[89]) | (~x[86] & x[87] & ~x[88] & ~x[89]) | (~x[86] & ~x[87] & x[88] & ~x[89]) | (~x[86] & ~x[87] & ~x[88] & x[89]) | (x[86] & x[87] & x[88] & ~x[89]) | (x[86] & x[87] & ~x[88] & x[89]) | (x[86] & ~x[87] & x[88] & x[89]) | (~x[86] & x[87] & x[88] & x[89]);
  assign t[323] = (x[87]);
  assign t[324] = (x[33]);
  assign t[325] = (x[62]);
  assign t[326] = (x[59]);
  assign t[327] = (x[68]);
  assign t[328] = (x[65]);
  assign t[329] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[32] = t[49] ^ t[31];
  assign t[330] = (x[98]);
  assign t[331] = (x[76]);
  assign t[332] = (x[73]);
  assign t[333] = (x[43]);
  assign t[334] = (x[51]);
  assign t[335] = (x[89]);
  assign t[336] = (x[86]);
  assign t[337] = (x[61]);
  assign t[338] = (x[67]);
  assign t[339] = (x[100]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[97]);
  assign t[341] = (x[75]);
  assign t[342] = (x[88]);
  assign t[343] = (x[99]);
  assign t[34] = t[52] ^ t[53];
  assign t[35] = ~(t[54] & t[55]);
  assign t[36] = ~(t[56] & t[117]);
  assign t[37] = t[57] ? x[38] : x[37];
  assign t[38] = ~(t[58] & t[59]);
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = t[66] ^ t[41];
  assign t[43] = ~(t[118]);
  assign t[44] = ~(t[119]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = ~(t[69]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[120]);
  assign t[49] = t[46] ? x[48] : x[47];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[121]);
  assign t[52] = t[46] ? x[56] : x[55];
  assign t[53] = ~(t[76] & t[77]);
  assign t[54] = ~(t[122]);
  assign t[55] = ~(t[123]);
  assign t[56] = ~(t[78] & t[79]);
  assign t[57] = ~(t[69]);
  assign t[58] = ~(t[80] & t[81]);
  assign t[59] = ~(t[82] & t[124]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[125]);
  assign t[62] = t[112] ? x[72] : x[71];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[126]);
  assign t[66] = t[112] ? x[80] : x[79];
  assign t[67] = ~(t[119] & t[118]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[112]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[91] & t[92]);
  assign t[73] = ~(t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[93] & t[94]);
  assign t[76] = ~(t[95] & t[96]);
  assign t[77] = ~(t[97] & t[132]);
  assign t[78] = ~(t[123] & t[122]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[98] & t[99]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[103]);
  assign t[87] = ~(t[104] & t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[140]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[105] & t[106]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[131] & t[130]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[144]);
  assign t[97] = ~(t[107] & t[108]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [106:0] x;
 output y;

 wire [277:0] t;
  assign t[0] = t[1] ? t[2] : t[90];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = t[154] ^ x[5];
  assign t[123] = t[155] ^ x[11];
  assign t[124] = t[156] ^ x[14];
  assign t[125] = t[157] ^ x[17];
  assign t[126] = t[158] ^ x[20];
  assign t[127] = t[159] ^ x[28];
  assign t[128] = t[160] ^ x[29];
  assign t[129] = t[161] ^ x[37];
  assign t[12] = t[93] ? x[21] : x[22];
  assign t[130] = t[162] ^ x[38];
  assign t[131] = t[163] ^ x[41];
  assign t[132] = t[164] ^ x[47];
  assign t[133] = t[165] ^ x[48];
  assign t[134] = t[166] ^ x[56];
  assign t[135] = t[167] ^ x[57];
  assign t[136] = t[168] ^ x[60];
  assign t[137] = t[169] ^ x[66];
  assign t[138] = t[170] ^ x[67];
  assign t[139] = t[171] ^ x[73];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = t[172] ^ x[74];
  assign t[141] = t[173] ^ x[82];
  assign t[142] = t[174] ^ x[83];
  assign t[143] = t[175] ^ x[86];
  assign t[144] = t[176] ^ x[92];
  assign t[145] = t[177] ^ x[93];
  assign t[146] = t[178] ^ x[94];
  assign t[147] = t[179] ^ x[95];
  assign t[148] = t[180] ^ x[96];
  assign t[149] = t[181] ^ x[97];
  assign t[14] = x[7] ? t[19] : t[18];
  assign t[150] = t[182] ^ x[103];
  assign t[151] = t[183] ^ x[104];
  assign t[152] = t[184] ^ x[105];
  assign t[153] = t[185] ^ x[106];
  assign t[154] = (~t[186] & t[187]);
  assign t[155] = (~t[188] & t[189]);
  assign t[156] = (~t[190] & t[191]);
  assign t[157] = (~t[192] & t[193]);
  assign t[158] = (~t[194] & t[195]);
  assign t[159] = (~t[196] & t[197]);
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = (~t[196] & t[198]);
  assign t[161] = (~t[199] & t[200]);
  assign t[162] = (~t[199] & t[201]);
  assign t[163] = (~t[196] & t[202]);
  assign t[164] = (~t[203] & t[204]);
  assign t[165] = (~t[203] & t[205]);
  assign t[166] = (~t[206] & t[207]);
  assign t[167] = (~t[206] & t[208]);
  assign t[168] = (~t[199] & t[209]);
  assign t[169] = (~t[210] & t[211]);
  assign t[16] = x[7] ? t[23] : t[22];
  assign t[170] = (~t[210] & t[212]);
  assign t[171] = (~t[213] & t[214]);
  assign t[172] = (~t[213] & t[215]);
  assign t[173] = (~t[216] & t[217]);
  assign t[174] = (~t[216] & t[218]);
  assign t[175] = (~t[203] & t[219]);
  assign t[176] = (~t[220] & t[221]);
  assign t[177] = (~t[220] & t[222]);
  assign t[178] = (~t[206] & t[223]);
  assign t[179] = (~t[210] & t[224]);
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = (~t[213] & t[225]);
  assign t[181] = (~t[216] & t[226]);
  assign t[182] = (~t[227] & t[228]);
  assign t[183] = (~t[227] & t[229]);
  assign t[184] = (~t[220] & t[230]);
  assign t[185] = (~t[227] & t[231]);
  assign t[186] = t[232] ^ x[4];
  assign t[187] = t[233] ^ x[5];
  assign t[188] = t[234] ^ x[10];
  assign t[189] = t[235] ^ x[11];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = t[236] ^ x[13];
  assign t[191] = t[237] ^ x[14];
  assign t[192] = t[238] ^ x[16];
  assign t[193] = t[239] ^ x[17];
  assign t[194] = t[240] ^ x[19];
  assign t[195] = t[241] ^ x[20];
  assign t[196] = t[242] ^ x[27];
  assign t[197] = t[243] ^ x[28];
  assign t[198] = t[244] ^ x[29];
  assign t[199] = t[245] ^ x[36];
  assign t[19] = t[28] ^ t[22];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[246] ^ x[37];
  assign t[201] = t[247] ^ x[38];
  assign t[202] = t[248] ^ x[41];
  assign t[203] = t[249] ^ x[46];
  assign t[204] = t[250] ^ x[47];
  assign t[205] = t[251] ^ x[48];
  assign t[206] = t[252] ^ x[55];
  assign t[207] = t[253] ^ x[56];
  assign t[208] = t[254] ^ x[57];
  assign t[209] = t[255] ^ x[60];
  assign t[20] = x[7] ? t[30] : t[29];
  assign t[210] = t[256] ^ x[65];
  assign t[211] = t[257] ^ x[66];
  assign t[212] = t[258] ^ x[67];
  assign t[213] = t[259] ^ x[72];
  assign t[214] = t[260] ^ x[73];
  assign t[215] = t[261] ^ x[74];
  assign t[216] = t[262] ^ x[81];
  assign t[217] = t[263] ^ x[82];
  assign t[218] = t[264] ^ x[83];
  assign t[219] = t[265] ^ x[86];
  assign t[21] = x[7] ? t[32] : t[31];
  assign t[220] = t[266] ^ x[91];
  assign t[221] = t[267] ^ x[92];
  assign t[222] = t[268] ^ x[93];
  assign t[223] = t[269] ^ x[94];
  assign t[224] = t[270] ^ x[95];
  assign t[225] = t[271] ^ x[96];
  assign t[226] = t[272] ^ x[97];
  assign t[227] = t[273] ^ x[102];
  assign t[228] = t[274] ^ x[103];
  assign t[229] = t[275] ^ x[104];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[276] ^ x[105];
  assign t[231] = t[277] ^ x[106];
  assign t[232] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[233] = (x[1]);
  assign t[234] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[235] = (x[9]);
  assign t[236] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[237] = (x[12]);
  assign t[238] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[239] = (x[15]);
  assign t[23] = t[35] ^ t[36];
  assign t[240] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[241] = (x[18]);
  assign t[242] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[243] = (x[25]);
  assign t[244] = (x[23]);
  assign t[245] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[246] = (x[34]);
  assign t[247] = (x[32]);
  assign t[248] = (x[26]);
  assign t[249] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = (x[44]);
  assign t[251] = (x[42]);
  assign t[252] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[253] = (x[53]);
  assign t[254] = (x[51]);
  assign t[255] = (x[35]);
  assign t[256] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[257] = (x[63]);
  assign t[258] = (x[61]);
  assign t[259] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = (x[70]);
  assign t[261] = (x[68]);
  assign t[262] = (x[77] & ~x[78] & ~x[79] & ~x[80]) | (~x[77] & x[78] & ~x[79] & ~x[80]) | (~x[77] & ~x[78] & x[79] & ~x[80]) | (~x[77] & ~x[78] & ~x[79] & x[80]) | (x[77] & x[78] & x[79] & ~x[80]) | (x[77] & x[78] & ~x[79] & x[80]) | (x[77] & ~x[78] & x[79] & x[80]) | (~x[77] & x[78] & x[79] & x[80]);
  assign t[263] = (x[79]);
  assign t[264] = (x[77]);
  assign t[265] = (x[45]);
  assign t[266] = (x[87] & ~x[88] & ~x[89] & ~x[90]) | (~x[87] & x[88] & ~x[89] & ~x[90]) | (~x[87] & ~x[88] & x[89] & ~x[90]) | (~x[87] & ~x[88] & ~x[89] & x[90]) | (x[87] & x[88] & x[89] & ~x[90]) | (x[87] & x[88] & ~x[89] & x[90]) | (x[87] & ~x[88] & x[89] & x[90]) | (~x[87] & x[88] & x[89] & x[90]);
  assign t[267] = (x[89]);
  assign t[268] = (x[87]);
  assign t[269] = (x[54]);
  assign t[26] = ~(t[95] & t[41]);
  assign t[270] = (x[64]);
  assign t[271] = (x[71]);
  assign t[272] = (x[80]);
  assign t[273] = (x[98] & ~x[99] & ~x[100] & ~x[101]) | (~x[98] & x[99] & ~x[100] & ~x[101]) | (~x[98] & ~x[99] & x[100] & ~x[101]) | (~x[98] & ~x[99] & ~x[100] & x[101]) | (x[98] & x[99] & x[100] & ~x[101]) | (x[98] & x[99] & ~x[100] & x[101]) | (x[98] & ~x[99] & x[100] & x[101]) | (~x[98] & x[99] & x[100] & x[101]);
  assign t[274] = (x[100]);
  assign t[275] = (x[98]);
  assign t[276] = (x[90]);
  assign t[277] = (x[101]);
  assign t[27] = ~(t[96] & t[42]);
  assign t[28] = t[43] ? x[31] : x[30];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[46] ^ t[47];
  assign t[31] = ~(t[48] & t[49]);
  assign t[32] = t[50] ^ t[31];
  assign t[33] = ~(t[97] & t[51]);
  assign t[34] = ~(t[98] & t[52]);
  assign t[35] = t[43] ? x[40] : x[39];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = ~(t[55] & t[56]);
  assign t[38] = t[57] ^ t[37];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[99]);
  assign t[42] = ~(t[99] & t[62]);
  assign t[43] = ~(t[63]);
  assign t[44] = ~(t[100] & t[64]);
  assign t[45] = ~(t[101] & t[65]);
  assign t[46] = t[43] ? x[50] : x[49];
  assign t[47] = ~(t[66] & t[67]);
  assign t[48] = ~(t[102] & t[68]);
  assign t[49] = ~(t[103] & t[69]);
  assign t[4] = ~(x[6]);
  assign t[50] = t[43] ? x[59] : x[58];
  assign t[51] = ~(t[104]);
  assign t[52] = ~(t[104] & t[70]);
  assign t[53] = ~(t[105] & t[71]);
  assign t[54] = ~(t[106] & t[72]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = ~(t[108] & t[74]);
  assign t[57] = t[93] ? x[76] : x[75];
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = ~(t[110] & t[76]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[93] ? x[85] : x[84];
  assign t[61] = ~(t[77] & t[78]);
  assign t[62] = ~(t[95]);
  assign t[63] = ~(t[93]);
  assign t[64] = ~(t[111]);
  assign t[65] = ~(t[111] & t[79]);
  assign t[66] = ~(t[112] & t[80]);
  assign t[67] = ~(t[113] & t[81]);
  assign t[68] = ~(t[114]);
  assign t[69] = ~(t[114] & t[82]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[97]);
  assign t[71] = ~(t[115]);
  assign t[72] = ~(t[115] & t[83]);
  assign t[73] = ~(t[116]);
  assign t[74] = ~(t[116] & t[84]);
  assign t[75] = ~(t[117]);
  assign t[76] = ~(t[117] & t[85]);
  assign t[77] = ~(t[118] & t[86]);
  assign t[78] = ~(t[119] & t[87]);
  assign t[79] = ~(t[100]);
  assign t[7] = ~(t[91] & t[92]);
  assign t[80] = ~(t[120]);
  assign t[81] = ~(t[120] & t[88]);
  assign t[82] = ~(t[102]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[107]);
  assign t[85] = ~(t[109]);
  assign t[86] = ~(t[121]);
  assign t[87] = ~(t[121] & t[89]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[118]);
  assign t[8] = ~(t[93] & t[94]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [115:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[223]);
  assign t[101] = ~(t[212] | t[213]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[142] | t[143]);
  assign t[105] = ~(t[144] | t[145]);
  assign t[106] = ~(t[226]);
  assign t[107] = ~(t[227]);
  assign t[108] = ~(t[146] | t[147]);
  assign t[109] = ~(t[148] | t[149]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[228] | t[150]);
  assign t[111] = t[151] ? x[100] : x[99];
  assign t[112] = ~(t[152] & t[153]);
  assign t[113] = ~(t[229]);
  assign t[114] = ~(t[230]);
  assign t[115] = ~(t[154] | t[155]);
  assign t[116] = t[204] ? x[104] : x[103];
  assign t[117] = t[156] | t[157];
  assign t[118] = ~(t[204]);
  assign t[119] = ~(t[158] & t[205]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[159] & t[160]);
  assign t[121] = ~(t[77] | t[161]);
  assign t[122] = ~(t[77] | t[162]);
  assign t[123] = t[205] & t[163];
  assign t[124] = t[159] | t[158];
  assign t[125] = ~(t[164] & t[160]);
  assign t[126] = ~(x[7] & t[165]);
  assign t[127] = ~(t[159] & t[205]);
  assign t[128] = ~(t[158] & t[160]);
  assign t[129] = ~(t[204]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[140]);
  assign t[131] = ~(t[231]);
  assign t[132] = ~(t[218] | t[219]);
  assign t[133] = ~(t[166] | t[144]);
  assign t[134] = ~(t[167] | t[168]);
  assign t[135] = ~(t[232]);
  assign t[136] = ~(t[220] | t[221]);
  assign t[137] = ~(t[233]);
  assign t[138] = ~(t[234]);
  assign t[139] = ~(t[169] | t[170]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[171] | t[144]);
  assign t[141] = ~(t[172] | t[173]);
  assign t[142] = ~(t[235]);
  assign t[143] = ~(t[224] | t[225]);
  assign t[144] = ~(t[118] | t[174]);
  assign t[145] = t[175] | t[176];
  assign t[146] = ~(t[236]);
  assign t[147] = ~(t[226] | t[227]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[238]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[177] | t[178]);
  assign t[151] = ~(t[129]);
  assign t[152] = ~(t[156] | t[179]);
  assign t[153] = ~(t[47]);
  assign t[154] = ~(t[239]);
  assign t[155] = ~(t[229] | t[230]);
  assign t[156] = ~(t[180] & t[181]);
  assign t[157] = ~(t[182] & t[86]);
  assign t[158] = x[7] & t[203];
  assign t[159] = ~(x[7] | t[203]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[205]);
  assign t[161] = t[202] ? t[119] : t[120];
  assign t[162] = t[202] ? t[184] : t[183];
  assign t[163] = ~(t[118] | t[202]);
  assign t[164] = ~(x[7] | t[185]);
  assign t[165] = ~(t[203] | t[160]);
  assign t[166] = ~(t[118] | t[186]);
  assign t[167] = ~(t[31]);
  assign t[168] = ~(t[77] | t[187]);
  assign t[169] = ~(t[240]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[233] | t[234]);
  assign t[171] = ~(t[118] | t[188]);
  assign t[172] = ~(t[189] & t[190]);
  assign t[173] = ~(t[80] & t[191]);
  assign t[174] = t[202] ? t[125] : t[184];
  assign t[175] = ~(t[77] | t[192]);
  assign t[176] = ~(t[180]);
  assign t[177] = ~(t[241]);
  assign t[178] = ~(t[237] | t[238]);
  assign t[179] = ~(t[193] & t[191]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[163] & t[194]);
  assign t[181] = ~(t[165] & t[195]);
  assign t[182] = ~(t[47] | t[175]);
  assign t[183] = ~(t[205] & t[164]);
  assign t[184] = ~(x[7] & t[196]);
  assign t[185] = ~(t[203]);
  assign t[186] = t[202] ? t[120] : t[128];
  assign t[187] = t[202] ? t[183] : t[184];
  assign t[188] = t[202] ? t[128] : t[120];
  assign t[189] = ~(t[166] | t[197]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[118] & t[198]);
  assign t[191] = t[118] | t[199];
  assign t[192] = t[202] ? t[127] : t[128];
  assign t[193] = ~(t[144]);
  assign t[194] = ~(t[183] & t[126]);
  assign t[195] = t[77] & t[202];
  assign t[196] = ~(t[203] | t[205]);
  assign t[197] = ~(t[77] | t[200]);
  assign t[198] = ~(t[184] & t[183]);
  assign t[199] = t[202] ? t[184] : t[125];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[125] : t[126];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[204] ? x[9] : x[10];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[32] | t[33]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[26] ^ t[34]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[5];
  assign t[243] = t[284] ^ x[13];
  assign t[244] = t[285] ^ x[16];
  assign t[245] = t[286] ^ x[19];
  assign t[246] = t[287] ^ x[22];
  assign t[247] = t[288] ^ x[28];
  assign t[248] = t[289] ^ x[34];
  assign t[249] = t[290] ^ x[35];
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = t[291] ^ x[36];
  assign t[251] = t[292] ^ x[44];
  assign t[252] = t[293] ^ x[50];
  assign t[253] = t[294] ^ x[51];
  assign t[254] = t[295] ^ x[52];
  assign t[255] = t[296] ^ x[58];
  assign t[256] = t[297] ^ x[66];
  assign t[257] = t[298] ^ x[72];
  assign t[258] = t[299] ^ x[73];
  assign t[259] = t[300] ^ x[74];
  assign t[25] = x[7] ? t[38] : t[37];
  assign t[260] = t[301] ^ x[75];
  assign t[261] = t[302] ^ x[78];
  assign t[262] = t[303] ^ x[79];
  assign t[263] = t[304] ^ x[85];
  assign t[264] = t[305] ^ x[88];
  assign t[265] = t[306] ^ x[89];
  assign t[266] = t[307] ^ x[90];
  assign t[267] = t[308] ^ x[91];
  assign t[268] = t[309] ^ x[92];
  assign t[269] = t[310] ^ x[98];
  assign t[26] = ~(t[39] | t[40]);
  assign t[270] = t[311] ^ x[101];
  assign t[271] = t[312] ^ x[102];
  assign t[272] = t[313] ^ x[105];
  assign t[273] = t[314] ^ x[106];
  assign t[274] = t[315] ^ x[107];
  assign t[275] = t[316] ^ x[108];
  assign t[276] = t[317] ^ x[109];
  assign t[277] = t[318] ^ x[110];
  assign t[278] = t[319] ^ x[111];
  assign t[279] = t[320] ^ x[112];
  assign t[27] = ~(t[41] ^ t[42]);
  assign t[280] = t[321] ^ x[113];
  assign t[281] = t[322] ^ x[114];
  assign t[282] = t[323] ^ x[115];
  assign t[283] = (~t[324] & t[325]);
  assign t[284] = (~t[326] & t[327]);
  assign t[285] = (~t[328] & t[329]);
  assign t[286] = (~t[330] & t[331]);
  assign t[287] = (~t[332] & t[333]);
  assign t[288] = (~t[334] & t[335]);
  assign t[289] = (~t[336] & t[337]);
  assign t[28] = x[7] ? t[44] : t[43];
  assign t[290] = (~t[334] & t[338]);
  assign t[291] = (~t[334] & t[339]);
  assign t[292] = (~t[340] & t[341]);
  assign t[293] = (~t[342] & t[343]);
  assign t[294] = (~t[336] & t[344]);
  assign t[295] = (~t[336] & t[345]);
  assign t[296] = (~t[346] & t[347]);
  assign t[297] = (~t[348] & t[349]);
  assign t[298] = (~t[350] & t[351]);
  assign t[299] = (~t[334] & t[352]);
  assign t[29] = x[7] ? t[46] : t[45];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[340] & t[353]);
  assign t[301] = (~t[340] & t[354]);
  assign t[302] = (~t[342] & t[355]);
  assign t[303] = (~t[342] & t[356]);
  assign t[304] = (~t[357] & t[358]);
  assign t[305] = (~t[336] & t[359]);
  assign t[306] = (~t[346] & t[360]);
  assign t[307] = (~t[346] & t[361]);
  assign t[308] = (~t[348] & t[362]);
  assign t[309] = (~t[348] & t[363]);
  assign t[30] = ~(t[47] | t[48]);
  assign t[310] = (~t[364] & t[365]);
  assign t[311] = (~t[350] & t[366]);
  assign t[312] = (~t[350] & t[367]);
  assign t[313] = (~t[340] & t[368]);
  assign t[314] = (~t[342] & t[369]);
  assign t[315] = (~t[357] & t[370]);
  assign t[316] = (~t[357] & t[371]);
  assign t[317] = (~t[346] & t[372]);
  assign t[318] = (~t[348] & t[373]);
  assign t[319] = (~t[364] & t[374]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (~t[364] & t[375]);
  assign t[321] = (~t[350] & t[376]);
  assign t[322] = (~t[357] & t[377]);
  assign t[323] = (~t[364] & t[378]);
  assign t[324] = t[379] ^ x[4];
  assign t[325] = t[380] ^ x[5];
  assign t[326] = t[381] ^ x[12];
  assign t[327] = t[382] ^ x[13];
  assign t[328] = t[383] ^ x[15];
  assign t[329] = t[384] ^ x[16];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[385] ^ x[18];
  assign t[331] = t[386] ^ x[19];
  assign t[332] = t[387] ^ x[21];
  assign t[333] = t[388] ^ x[22];
  assign t[334] = t[389] ^ x[27];
  assign t[335] = t[390] ^ x[28];
  assign t[336] = t[391] ^ x[33];
  assign t[337] = t[392] ^ x[34];
  assign t[338] = t[393] ^ x[35];
  assign t[339] = t[394] ^ x[36];
  assign t[33] = ~(t[206] | t[53]);
  assign t[340] = t[395] ^ x[43];
  assign t[341] = t[396] ^ x[44];
  assign t[342] = t[397] ^ x[49];
  assign t[343] = t[398] ^ x[50];
  assign t[344] = t[399] ^ x[51];
  assign t[345] = t[400] ^ x[52];
  assign t[346] = t[401] ^ x[57];
  assign t[347] = t[402] ^ x[58];
  assign t[348] = t[403] ^ x[65];
  assign t[349] = t[404] ^ x[66];
  assign t[34] = ~(t[54] ^ t[55]);
  assign t[350] = t[405] ^ x[71];
  assign t[351] = t[406] ^ x[72];
  assign t[352] = t[407] ^ x[73];
  assign t[353] = t[408] ^ x[74];
  assign t[354] = t[409] ^ x[75];
  assign t[355] = t[410] ^ x[78];
  assign t[356] = t[411] ^ x[79];
  assign t[357] = t[412] ^ x[84];
  assign t[358] = t[413] ^ x[85];
  assign t[359] = t[414] ^ x[88];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[415] ^ x[89];
  assign t[361] = t[416] ^ x[90];
  assign t[362] = t[417] ^ x[91];
  assign t[363] = t[418] ^ x[92];
  assign t[364] = t[419] ^ x[97];
  assign t[365] = t[420] ^ x[98];
  assign t[366] = t[421] ^ x[101];
  assign t[367] = t[422] ^ x[102];
  assign t[368] = t[423] ^ x[105];
  assign t[369] = t[424] ^ x[106];
  assign t[36] = ~(t[35] ^ t[58]);
  assign t[370] = t[425] ^ x[107];
  assign t[371] = t[426] ^ x[108];
  assign t[372] = t[427] ^ x[109];
  assign t[373] = t[428] ^ x[110];
  assign t[374] = t[429] ^ x[111];
  assign t[375] = t[430] ^ x[112];
  assign t[376] = t[431] ^ x[113];
  assign t[377] = t[432] ^ x[114];
  assign t[378] = t[433] ^ x[115];
  assign t[379] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = ~(t[59] | t[60]);
  assign t[380] = (x[0]);
  assign t[381] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[382] = (x[11]);
  assign t[383] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[384] = (x[14]);
  assign t[385] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[386] = (x[17]);
  assign t[387] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[388] = (x[20]);
  assign t[389] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[38] = ~(t[61] ^ t[62]);
  assign t[390] = (x[24]);
  assign t[391] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[392] = (x[30]);
  assign t[393] = (x[25]);
  assign t[394] = (x[26]);
  assign t[395] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[396] = (x[40]);
  assign t[397] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[398] = (x[46]);
  assign t[399] = (x[31]);
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[32]);
  assign t[401] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[402] = (x[54]);
  assign t[403] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[404] = (x[62]);
  assign t[405] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[406] = (x[68]);
  assign t[407] = (x[23]);
  assign t[408] = (x[41]);
  assign t[409] = (x[42]);
  assign t[40] = ~(t[207] | t[65]);
  assign t[410] = (x[47]);
  assign t[411] = (x[48]);
  assign t[412] = (x[80] & ~x[81] & ~x[82] & ~x[83]) | (~x[80] & x[81] & ~x[82] & ~x[83]) | (~x[80] & ~x[81] & x[82] & ~x[83]) | (~x[80] & ~x[81] & ~x[82] & x[83]) | (x[80] & x[81] & x[82] & ~x[83]) | (x[80] & x[81] & ~x[82] & x[83]) | (x[80] & ~x[81] & x[82] & x[83]) | (~x[80] & x[81] & x[82] & x[83]);
  assign t[413] = (x[81]);
  assign t[414] = (x[29]);
  assign t[415] = (x[55]);
  assign t[416] = (x[56]);
  assign t[417] = (x[63]);
  assign t[418] = (x[64]);
  assign t[419] = (x[93] & ~x[94] & ~x[95] & ~x[96]) | (~x[93] & x[94] & ~x[95] & ~x[96]) | (~x[93] & ~x[94] & x[95] & ~x[96]) | (~x[93] & ~x[94] & ~x[95] & x[96]) | (x[93] & x[94] & x[95] & ~x[96]) | (x[93] & x[94] & ~x[95] & x[96]) | (x[93] & ~x[94] & x[95] & x[96]) | (~x[93] & x[94] & x[95] & x[96]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (x[94]);
  assign t[421] = (x[69]);
  assign t[422] = (x[70]);
  assign t[423] = (x[39]);
  assign t[424] = (x[45]);
  assign t[425] = (x[82]);
  assign t[426] = (x[83]);
  assign t[427] = (x[53]);
  assign t[428] = (x[61]);
  assign t[429] = (x[95]);
  assign t[42] = ~(t[68] ^ t[69]);
  assign t[430] = (x[96]);
  assign t[431] = (x[67]);
  assign t[432] = (x[80]);
  assign t[433] = (x[93]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[46] = ~(t[45] ^ t[76]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[48] = ~(t[79] & t[80]);
  assign t[49] = ~(t[77] | t[81]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[77] | t[82]);
  assign t[51] = ~(t[208]);
  assign t[52] = ~(t[209]);
  assign t[53] = ~(t[83] | t[84]);
  assign t[54] = t[85] ? x[38] : x[37];
  assign t[55] = ~(t[86] & t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[210] | t[90]);
  assign t[58] = ~(t[91] ^ t[92]);
  assign t[59] = ~(t[93] | t[94]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[211] | t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[212]);
  assign t[64] = ~(t[213]);
  assign t[65] = ~(t[100] | t[101]);
  assign t[66] = ~(t[102] | t[103]);
  assign t[67] = ~(t[214] | t[104]);
  assign t[68] = t[204] ? x[60] : x[59];
  assign t[69] = ~(t[30] & t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[215] | t[108]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[111] ^ t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[216] | t[115]);
  assign t[76] = ~(t[116] ^ t[117]);
  assign t[77] = ~(t[118]);
  assign t[78] = t[202] ? t[120] : t[119];
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[123] & t[124]);
  assign t[81] = t[202] ? t[126] : t[125];
  assign t[82] = t[202] ? t[128] : t[127];
  assign t[83] = ~(t[217]);
  assign t[84] = ~(t[208] | t[209]);
  assign t[85] = ~(t[129]);
  assign t[86] = ~(t[122] | t[50]);
  assign t[87] = ~(t[123] | t[130]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[219]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = t[85] ? x[77] : x[76];
  assign t[92] = ~(t[133] & t[134]);
  assign t[93] = ~(t[220]);
  assign t[94] = ~(t[221]);
  assign t[95] = ~(t[135] | t[136]);
  assign t[96] = ~(t[137] | t[138]);
  assign t[97] = ~(t[222] | t[139]);
  assign t[98] = t[85] ? x[87] : x[86];
  assign t[99] = ~(t[140] & t[141]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [172:0] x;
 output y;

 wire [672:0] t;
  assign t[0] = t[1] ? t[2] : t[403];
  assign t[100] = ~(t[425] | t[145]);
  assign t[101] = t[146] ? x[91] : x[90];
  assign t[102] = ~(t[147] & t[83]);
  assign t[103] = ~(t[426]);
  assign t[104] = ~(t[427]);
  assign t[105] = ~(t[148] | t[149]);
  assign t[106] = t[146] ? x[95] : x[94];
  assign t[107] = ~(t[150] & t[151]);
  assign t[108] = ~(t[428]);
  assign t[109] = ~(t[415] | t[416]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[429]);
  assign t[111] = ~(t[430]);
  assign t[112] = ~(t[152] | t[153]);
  assign t[113] = ~(t[154] | t[155]);
  assign t[114] = ~(t[431]);
  assign t[115] = ~(t[432]);
  assign t[116] = ~(t[156] | t[157]);
  assign t[117] = ~(t[158] | t[159]);
  assign t[118] = ~(t[433] | t[160]);
  assign t[119] = t[93] ? x[108] : x[107];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[161] & t[162]);
  assign t[121] = ~(t[434]);
  assign t[122] = ~(t[435]);
  assign t[123] = ~(t[163] | t[164]);
  assign t[124] = t[406] ? x[112] : x[111];
  assign t[125] = t[165] | t[166];
  assign t[126] = ~(t[167] & t[407]);
  assign t[127] = ~(t[168] & t[169]);
  assign t[128] = ~(t[80] | t[170]);
  assign t[129] = ~(t[80] | t[171]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[407] & t[172];
  assign t[131] = t[168] | t[167];
  assign t[132] = ~(x[7] & t[173]);
  assign t[133] = ~(t[174] & t[169]);
  assign t[134] = t[404] ? t[176] : t[175];
  assign t[135] = ~(t[172] & t[177]);
  assign t[136] = ~(t[436]);
  assign t[137] = ~(t[421] | t[422]);
  assign t[138] = ~(t[406]);
  assign t[139] = ~(t[113]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[80] | t[178]);
  assign t[141] = ~(t[437]);
  assign t[142] = ~(t[423] | t[424]);
  assign t[143] = ~(t[438]);
  assign t[144] = ~(t[439]);
  assign t[145] = ~(t[179] | t[180]);
  assign t[146] = ~(t[138]);
  assign t[147] = ~(t[165] | t[181]);
  assign t[148] = ~(t[440]);
  assign t[149] = ~(t[426] | t[427]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[128] | t[182]);
  assign t[151] = ~(t[183] & t[184]);
  assign t[152] = ~(t[441]);
  assign t[153] = ~(t[429] | t[430]);
  assign t[154] = ~(t[80] | t[185]);
  assign t[155] = ~(t[80] | t[186]);
  assign t[156] = ~(t[442]);
  assign t[157] = ~(t[431] | t[432]);
  assign t[158] = ~(t[443]);
  assign t[159] = ~(t[444]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[187] | t[188]);
  assign t[161] = ~(t[165] | t[189]);
  assign t[162] = ~(t[48]);
  assign t[163] = ~(t[445]);
  assign t[164] = ~(t[434] | t[435]);
  assign t[165] = ~(t[135] & t[151]);
  assign t[166] = ~(t[190] & t[191]);
  assign t[167] = x[7] & t[405];
  assign t[168] = ~(x[7] | t[405]);
  assign t[169] = ~(t[407]);
  assign t[16] = ~(t[404] & t[405]);
  assign t[170] = t[404] ? t[126] : t[127];
  assign t[171] = t[404] ? t[132] : t[192];
  assign t[172] = ~(t[84] | t[404]);
  assign t[173] = ~(t[405] | t[407]);
  assign t[174] = ~(x[7] | t[193]);
  assign t[175] = ~(t[167] & t[169]);
  assign t[176] = ~(t[168] & t[407]);
  assign t[177] = ~(t[192] & t[194]);
  assign t[178] = t[404] ? t[192] : t[132];
  assign t[179] = ~(t[446]);
  assign t[17] = ~(t[406] & t[407]);
  assign t[180] = ~(t[438] | t[439]);
  assign t[181] = t[140] | t[86];
  assign t[182] = ~(t[195] & t[196]);
  assign t[183] = ~(t[405] | t[169]);
  assign t[184] = t[80] & t[404];
  assign t[185] = t[404] ? t[194] : t[133];
  assign t[186] = t[404] ? t[175] : t[176];
  assign t[187] = ~(t[447]);
  assign t[188] = ~(t[443] | t[444]);
  assign t[189] = ~(t[197] & t[198]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[48] | t[86]);
  assign t[191] = ~(t[129] | t[155]);
  assign t[192] = ~(t[407] & t[174]);
  assign t[193] = ~(t[405]);
  assign t[194] = ~(x[7] & t[183]);
  assign t[195] = ~(t[199] | t[200]);
  assign t[196] = ~(t[84] & t[201]);
  assign t[197] = ~(t[50]);
  assign t[198] = t[84] | t[202];
  assign t[199] = ~(t[84] | t[203]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[80] | t[204]);
  assign t[201] = ~(t[132] & t[192]);
  assign t[202] = t[404] ? t[132] : t[133];
  assign t[203] = t[404] ? t[127] : t[175];
  assign t[204] = t[404] ? t[133] : t[194];
  assign t[205] = t[6] ? t[206] : t[448];
  assign t[206] = x[6] ? t[208] : t[207];
  assign t[207] = x[7] ? t[210] : t[209];
  assign t[208] = t[211] ^ x[126];
  assign t[209] = t[212] ^ t[213];
  assign t[20] = t[406] ? x[9] : x[10];
  assign t[210] = ~(t[214] ^ t[215]);
  assign t[211] = x[127] ^ x[128];
  assign t[212] = t[216] ? x[127] : x[128];
  assign t[213] = ~(t[217] ^ t[218]);
  assign t[214] = x[7] ? t[220] : t[219];
  assign t[215] = ~(t[221] ^ t[222]);
  assign t[216] = ~(t[138]);
  assign t[217] = x[7] ? t[224] : t[223];
  assign t[218] = ~(t[225] ^ t[226]);
  assign t[219] = ~(t[227] & t[228]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[229] ^ t[230];
  assign t[221] = x[7] ? t[232] : t[231];
  assign t[222] = x[7] ? t[234] : t[233];
  assign t[223] = ~(t[235] & t[236]);
  assign t[224] = t[237] ^ t[238];
  assign t[225] = x[7] ? t[240] : t[239];
  assign t[226] = x[7] ? t[242] : t[241];
  assign t[227] = ~(t[410] & t[53]);
  assign t[228] = ~(t[420] & t[243]);
  assign t[229] = t[93] ? x[130] : x[129];
  assign t[22] = ~(t[32] | t[33]);
  assign t[230] = ~(t[244] & t[245]);
  assign t[231] = ~(t[246] & t[247]);
  assign t[232] = t[248] ^ t[241];
  assign t[233] = ~(t[249] & t[250]);
  assign t[234] = t[251] ^ t[252];
  assign t[235] = ~(t[415] & t[67]);
  assign t[236] = ~(t[428] & t[253]);
  assign t[237] = t[406] ? x[132] : x[131];
  assign t[238] = ~(t[254] & t[255]);
  assign t[239] = ~(t[256] & t[257]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = t[258] ^ t[239];
  assign t[241] = ~(t[259] & t[260]);
  assign t[242] = t[261] ^ t[262];
  assign t[243] = ~(t[411] & t[52]);
  assign t[244] = ~(t[421] & t[91]);
  assign t[245] = ~(t[436] & t[263]);
  assign t[246] = ~(t[426] & t[104]);
  assign t[247] = ~(t[440] & t[264]);
  assign t[248] = t[146] ? x[134] : x[133];
  assign t[249] = ~(t[423] & t[97]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = ~(t[437] & t[265]);
  assign t[251] = t[146] ? x[136] : x[135];
  assign t[252] = ~(t[266] & t[267]);
  assign t[253] = ~(t[416] & t[66]);
  assign t[254] = ~(t[429] & t[111]);
  assign t[255] = ~(t[441] & t[268]);
  assign t[256] = ~(t[434] & t[122]);
  assign t[257] = ~(t[445] & t[269]);
  assign t[258] = t[406] ? x[138] : x[137];
  assign t[259] = ~(t[431] & t[115]);
  assign t[25] = x[7] ? t[39] : t[38];
  assign t[260] = ~(t[442] & t[270]);
  assign t[261] = t[406] ? x[140] : x[139];
  assign t[262] = ~(t[271] & t[272]);
  assign t[263] = ~(t[422] & t[90]);
  assign t[264] = ~(t[427] & t[103]);
  assign t[265] = ~(t[424] & t[96]);
  assign t[266] = ~(t[438] & t[144]);
  assign t[267] = ~(t[446] & t[273]);
  assign t[268] = ~(t[430] & t[110]);
  assign t[269] = ~(t[435] & t[121]);
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = ~(t[432] & t[114]);
  assign t[271] = ~(t[443] & t[159]);
  assign t[272] = ~(t[447] & t[274]);
  assign t[273] = ~(t[439] & t[143]);
  assign t[274] = ~(t[444] & t[158]);
  assign t[275] = t[6] ? t[276] : t[449];
  assign t[276] = x[6] ? t[278] : t[277];
  assign t[277] = x[7] ? t[280] : t[279];
  assign t[278] = t[281] ^ x[142];
  assign t[279] = t[282] ^ t[283];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = ~(t[284] ^ t[285]);
  assign t[281] = x[143] ^ x[144];
  assign t[282] = t[146] ? x[143] : x[144];
  assign t[283] = ~(t[286] ^ t[287]);
  assign t[284] = x[7] ? t[289] : t[288];
  assign t[285] = ~(t[290] ^ t[291]);
  assign t[286] = x[7] ? t[293] : t[292];
  assign t[287] = ~(t[294] ^ t[295]);
  assign t[288] = ~(t[296] & t[297]);
  assign t[289] = t[298] ^ t[299];
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = x[7] ? t[301] : t[300];
  assign t[291] = x[7] ? t[303] : t[302];
  assign t[292] = ~(t[304] & t[305]);
  assign t[293] = t[306] ^ t[307];
  assign t[294] = x[7] ? t[309] : t[308];
  assign t[295] = x[7] ? t[311] : t[310];
  assign t[296] = ~(t[53] & t[88]);
  assign t[297] = ~(t[312] & t[408]);
  assign t[298] = t[93] ? x[146] : x[145];
  assign t[299] = ~(t[313] & t[314]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = ~(t[315] & t[316]);
  assign t[301] = t[317] ^ t[308];
  assign t[302] = ~(t[318] & t[319]);
  assign t[303] = t[320] ^ t[321];
  assign t[304] = ~(t[67] & t[108]);
  assign t[305] = ~(t[322] & t[409]);
  assign t[306] = t[406] ? x[148] : x[147];
  assign t[307] = ~(t[323] & t[324]);
  assign t[308] = ~(t[325] & t[326]);
  assign t[309] = t[327] ^ t[328];
  assign t[30] = ~(t[48] | t[49]);
  assign t[310] = ~(t[329] & t[330]);
  assign t[311] = t[331] ^ t[310];
  assign t[312] = ~(t[332] & t[52]);
  assign t[313] = ~(t[91] & t[136]);
  assign t[314] = ~(t[333] & t[412]);
  assign t[315] = ~(t[104] & t[148]);
  assign t[316] = ~(t[334] & t[414]);
  assign t[317] = t[146] ? x[150] : x[149];
  assign t[318] = ~(t[97] & t[141]);
  assign t[319] = ~(t[335] & t[413]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = t[146] ? x[152] : x[151];
  assign t[321] = ~(t[336] & t[337]);
  assign t[322] = ~(t[338] & t[66]);
  assign t[323] = ~(t[111] & t[152]);
  assign t[324] = ~(t[339] & t[417]);
  assign t[325] = ~(t[115] & t[156]);
  assign t[326] = ~(t[340] & t[418]);
  assign t[327] = t[406] ? x[154] : x[153];
  assign t[328] = ~(t[341] & t[342]);
  assign t[329] = ~(t[122] & t[163]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = ~(t[343] & t[419]);
  assign t[331] = t[406] ? x[156] : x[155];
  assign t[332] = ~(t[420] & t[411]);
  assign t[333] = ~(t[344] & t[90]);
  assign t[334] = ~(t[345] & t[103]);
  assign t[335] = ~(t[346] & t[96]);
  assign t[336] = ~(t[144] & t[179]);
  assign t[337] = ~(t[347] & t[425]);
  assign t[338] = ~(t[428] & t[416]);
  assign t[339] = ~(t[348] & t[110]);
  assign t[33] = ~(t[408] | t[54]);
  assign t[340] = ~(t[349] & t[114]);
  assign t[341] = ~(t[159] & t[187]);
  assign t[342] = ~(t[350] & t[433]);
  assign t[343] = ~(t[351] & t[121]);
  assign t[344] = ~(t[436] & t[422]);
  assign t[345] = ~(t[440] & t[427]);
  assign t[346] = ~(t[437] & t[424]);
  assign t[347] = ~(t[352] & t[143]);
  assign t[348] = ~(t[441] & t[430]);
  assign t[349] = ~(t[442] & t[432]);
  assign t[34] = ~(t[55] | t[56]);
  assign t[350] = ~(t[353] & t[158]);
  assign t[351] = ~(t[445] & t[435]);
  assign t[352] = ~(t[446] & t[439]);
  assign t[353] = ~(t[447] & t[444]);
  assign t[354] = t[6] ? t[355] : t[450];
  assign t[355] = x[6] ? t[357] : t[356];
  assign t[356] = x[7] ? t[359] : t[358];
  assign t[357] = t[360] ^ x[158];
  assign t[358] = t[361] ^ t[362];
  assign t[359] = ~(t[363] ^ t[364]);
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[360] = x[159] ^ x[160];
  assign t[361] = t[93] ? x[160] : x[159];
  assign t[362] = ~(t[365] ^ t[366]);
  assign t[363] = x[7] ? t[368] : t[367];
  assign t[364] = ~(t[369] ^ t[370]);
  assign t[365] = x[7] ? t[372] : t[371];
  assign t[366] = ~(t[373] ^ t[374]);
  assign t[367] = ~(t[296] & t[375]);
  assign t[368] = t[376] ^ t[377];
  assign t[369] = x[7] ? t[379] : t[378];
  assign t[36] = ~(t[59] | t[60]);
  assign t[370] = x[7] ? t[381] : t[380];
  assign t[371] = ~(t[304] & t[382]);
  assign t[372] = t[383] ^ t[384];
  assign t[373] = x[7] ? t[386] : t[385];
  assign t[374] = x[7] ? t[388] : t[387];
  assign t[375] = t[32] | t[408];
  assign t[376] = t[93] ? x[162] : x[161];
  assign t[377] = ~(t[313] & t[389]);
  assign t[378] = ~(t[315] & t[390]);
  assign t[379] = t[391] ^ t[385];
  assign t[37] = ~(t[61] ^ t[62]);
  assign t[380] = ~(t[318] & t[392]);
  assign t[381] = t[393] ^ t[394];
  assign t[382] = t[40] | t[409];
  assign t[383] = t[406] ? x[164] : x[163];
  assign t[384] = ~(t[323] & t[395]);
  assign t[385] = ~(t[325] & t[396]);
  assign t[386] = t[397] ^ t[398];
  assign t[387] = ~(t[329] & t[399]);
  assign t[388] = t[400] ^ t[387];
  assign t[389] = t[55] | t[412];
  assign t[38] = ~(t[63] | t[64]);
  assign t[390] = t[63] | t[414];
  assign t[391] = t[146] ? x[166] : x[165];
  assign t[392] = t[59] | t[413];
  assign t[393] = t[146] ? x[168] : x[167];
  assign t[394] = ~(t[336] & t[401]);
  assign t[395] = t[69] | t[417];
  assign t[396] = t[73] | t[418];
  assign t[397] = t[406] ? x[170] : x[169];
  assign t[398] = ~(t[341] & t[402]);
  assign t[399] = t[77] | t[419];
  assign t[39] = ~(t[44] ^ t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[406] ? x[172] : x[171];
  assign t[401] = t[99] | t[425];
  assign t[402] = t[117] | t[433];
  assign t[403] = (t[451]);
  assign t[404] = (t[452]);
  assign t[405] = (t[453]);
  assign t[406] = (t[454]);
  assign t[407] = (t[455]);
  assign t[408] = (t[456]);
  assign t[409] = (t[457]);
  assign t[40] = ~(t[66] | t[67]);
  assign t[410] = (t[458]);
  assign t[411] = (t[459]);
  assign t[412] = (t[460]);
  assign t[413] = (t[461]);
  assign t[414] = (t[462]);
  assign t[415] = (t[463]);
  assign t[416] = (t[464]);
  assign t[417] = (t[465]);
  assign t[418] = (t[466]);
  assign t[419] = (t[467]);
  assign t[41] = ~(t[409] | t[68]);
  assign t[420] = (t[468]);
  assign t[421] = (t[469]);
  assign t[422] = (t[470]);
  assign t[423] = (t[471]);
  assign t[424] = (t[472]);
  assign t[425] = (t[473]);
  assign t[426] = (t[474]);
  assign t[427] = (t[475]);
  assign t[428] = (t[476]);
  assign t[429] = (t[477]);
  assign t[42] = ~(t[69] | t[70]);
  assign t[430] = (t[478]);
  assign t[431] = (t[479]);
  assign t[432] = (t[480]);
  assign t[433] = (t[481]);
  assign t[434] = (t[482]);
  assign t[435] = (t[483]);
  assign t[436] = (t[484]);
  assign t[437] = (t[485]);
  assign t[438] = (t[486]);
  assign t[439] = (t[487]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[440] = (t[488]);
  assign t[441] = (t[489]);
  assign t[442] = (t[490]);
  assign t[443] = (t[491]);
  assign t[444] = (t[492]);
  assign t[445] = (t[493]);
  assign t[446] = (t[494]);
  assign t[447] = (t[495]);
  assign t[448] = (t[496]);
  assign t[449] = (t[497]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[450] = (t[498]);
  assign t[451] = t[499] ^ x[5];
  assign t[452] = t[500] ^ x[13];
  assign t[453] = t[501] ^ x[16];
  assign t[454] = t[502] ^ x[19];
  assign t[455] = t[503] ^ x[22];
  assign t[456] = t[504] ^ x[28];
  assign t[457] = t[505] ^ x[34];
  assign t[458] = t[506] ^ x[35];
  assign t[459] = t[507] ^ x[36];
  assign t[45] = ~(t[75] ^ t[76]);
  assign t[460] = t[508] ^ x[42];
  assign t[461] = t[509] ^ x[50];
  assign t[462] = t[510] ^ x[56];
  assign t[463] = t[511] ^ x[57];
  assign t[464] = t[512] ^ x[58];
  assign t[465] = t[513] ^ x[64];
  assign t[466] = t[514] ^ x[72];
  assign t[467] = t[515] ^ x[78];
  assign t[468] = t[516] ^ x[79];
  assign t[469] = t[517] ^ x[80];
  assign t[46] = ~(t[77] | t[78]);
  assign t[470] = t[518] ^ x[81];
  assign t[471] = t[519] ^ x[82];
  assign t[472] = t[520] ^ x[83];
  assign t[473] = t[521] ^ x[89];
  assign t[474] = t[522] ^ x[92];
  assign t[475] = t[523] ^ x[93];
  assign t[476] = t[524] ^ x[96];
  assign t[477] = t[525] ^ x[97];
  assign t[478] = t[526] ^ x[98];
  assign t[479] = t[527] ^ x[99];
  assign t[47] = ~(t[46] ^ t[79]);
  assign t[480] = t[528] ^ x[100];
  assign t[481] = t[529] ^ x[106];
  assign t[482] = t[530] ^ x[109];
  assign t[483] = t[531] ^ x[110];
  assign t[484] = t[532] ^ x[113];
  assign t[485] = t[533] ^ x[114];
  assign t[486] = t[534] ^ x[115];
  assign t[487] = t[535] ^ x[116];
  assign t[488] = t[536] ^ x[117];
  assign t[489] = t[537] ^ x[118];
  assign t[48] = ~(t[80] | t[81]);
  assign t[490] = t[538] ^ x[119];
  assign t[491] = t[539] ^ x[120];
  assign t[492] = t[540] ^ x[121];
  assign t[493] = t[541] ^ x[122];
  assign t[494] = t[542] ^ x[123];
  assign t[495] = t[543] ^ x[124];
  assign t[496] = t[544] ^ x[125];
  assign t[497] = t[545] ^ x[141];
  assign t[498] = t[546] ^ x[157];
  assign t[499] = (~t[547] & t[548]);
  assign t[49] = ~(t[82] & t[83]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[549] & t[550]);
  assign t[501] = (~t[551] & t[552]);
  assign t[502] = (~t[553] & t[554]);
  assign t[503] = (~t[555] & t[556]);
  assign t[504] = (~t[557] & t[558]);
  assign t[505] = (~t[559] & t[560]);
  assign t[506] = (~t[557] & t[561]);
  assign t[507] = (~t[557] & t[562]);
  assign t[508] = (~t[563] & t[564]);
  assign t[509] = (~t[565] & t[566]);
  assign t[50] = ~(t[84] | t[85]);
  assign t[510] = (~t[567] & t[568]);
  assign t[511] = (~t[559] & t[569]);
  assign t[512] = (~t[559] & t[570]);
  assign t[513] = (~t[571] & t[572]);
  assign t[514] = (~t[573] & t[574]);
  assign t[515] = (~t[575] & t[576]);
  assign t[516] = (~t[557] & t[577]);
  assign t[517] = (~t[563] & t[578]);
  assign t[518] = (~t[563] & t[579]);
  assign t[519] = (~t[565] & t[580]);
  assign t[51] = t[86] | t[87];
  assign t[520] = (~t[565] & t[581]);
  assign t[521] = (~t[582] & t[583]);
  assign t[522] = (~t[567] & t[584]);
  assign t[523] = (~t[567] & t[585]);
  assign t[524] = (~t[559] & t[586]);
  assign t[525] = (~t[571] & t[587]);
  assign t[526] = (~t[571] & t[588]);
  assign t[527] = (~t[573] & t[589]);
  assign t[528] = (~t[573] & t[590]);
  assign t[529] = (~t[591] & t[592]);
  assign t[52] = ~(t[410]);
  assign t[530] = (~t[575] & t[593]);
  assign t[531] = (~t[575] & t[594]);
  assign t[532] = (~t[563] & t[595]);
  assign t[533] = (~t[565] & t[596]);
  assign t[534] = (~t[582] & t[597]);
  assign t[535] = (~t[582] & t[598]);
  assign t[536] = (~t[567] & t[599]);
  assign t[537] = (~t[571] & t[600]);
  assign t[538] = (~t[573] & t[601]);
  assign t[539] = (~t[591] & t[602]);
  assign t[53] = ~(t[411]);
  assign t[540] = (~t[591] & t[603]);
  assign t[541] = (~t[575] & t[604]);
  assign t[542] = (~t[582] & t[605]);
  assign t[543] = (~t[591] & t[606]);
  assign t[544] = (~t[547] & t[607]);
  assign t[545] = (~t[547] & t[608]);
  assign t[546] = (~t[547] & t[609]);
  assign t[547] = t[610] ^ x[4];
  assign t[548] = t[611] ^ x[5];
  assign t[549] = t[612] ^ x[12];
  assign t[54] = ~(t[88] | t[89]);
  assign t[550] = t[613] ^ x[13];
  assign t[551] = t[614] ^ x[15];
  assign t[552] = t[615] ^ x[16];
  assign t[553] = t[616] ^ x[18];
  assign t[554] = t[617] ^ x[19];
  assign t[555] = t[618] ^ x[21];
  assign t[556] = t[619] ^ x[22];
  assign t[557] = t[620] ^ x[27];
  assign t[558] = t[621] ^ x[28];
  assign t[559] = t[622] ^ x[33];
  assign t[55] = ~(t[90] | t[91]);
  assign t[560] = t[623] ^ x[34];
  assign t[561] = t[624] ^ x[35];
  assign t[562] = t[625] ^ x[36];
  assign t[563] = t[626] ^ x[41];
  assign t[564] = t[627] ^ x[42];
  assign t[565] = t[628] ^ x[49];
  assign t[566] = t[629] ^ x[50];
  assign t[567] = t[630] ^ x[55];
  assign t[568] = t[631] ^ x[56];
  assign t[569] = t[632] ^ x[57];
  assign t[56] = ~(t[412] | t[92]);
  assign t[570] = t[633] ^ x[58];
  assign t[571] = t[634] ^ x[63];
  assign t[572] = t[635] ^ x[64];
  assign t[573] = t[636] ^ x[71];
  assign t[574] = t[637] ^ x[72];
  assign t[575] = t[638] ^ x[77];
  assign t[576] = t[639] ^ x[78];
  assign t[577] = t[640] ^ x[79];
  assign t[578] = t[641] ^ x[80];
  assign t[579] = t[642] ^ x[81];
  assign t[57] = t[93] ? x[44] : x[43];
  assign t[580] = t[643] ^ x[82];
  assign t[581] = t[644] ^ x[83];
  assign t[582] = t[645] ^ x[88];
  assign t[583] = t[646] ^ x[89];
  assign t[584] = t[647] ^ x[92];
  assign t[585] = t[648] ^ x[93];
  assign t[586] = t[649] ^ x[96];
  assign t[587] = t[650] ^ x[97];
  assign t[588] = t[651] ^ x[98];
  assign t[589] = t[652] ^ x[99];
  assign t[58] = ~(t[94] & t[95]);
  assign t[590] = t[653] ^ x[100];
  assign t[591] = t[654] ^ x[105];
  assign t[592] = t[655] ^ x[106];
  assign t[593] = t[656] ^ x[109];
  assign t[594] = t[657] ^ x[110];
  assign t[595] = t[658] ^ x[113];
  assign t[596] = t[659] ^ x[114];
  assign t[597] = t[660] ^ x[115];
  assign t[598] = t[661] ^ x[116];
  assign t[599] = t[662] ^ x[117];
  assign t[59] = ~(t[96] | t[97]);
  assign t[5] = t[9] ^ x[8];
  assign t[600] = t[663] ^ x[118];
  assign t[601] = t[664] ^ x[119];
  assign t[602] = t[665] ^ x[120];
  assign t[603] = t[666] ^ x[121];
  assign t[604] = t[667] ^ x[122];
  assign t[605] = t[668] ^ x[123];
  assign t[606] = t[669] ^ x[124];
  assign t[607] = t[670] ^ x[125];
  assign t[608] = t[671] ^ x[141];
  assign t[609] = t[672] ^ x[157];
  assign t[60] = ~(t[413] | t[98]);
  assign t[610] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[611] = (x[0]);
  assign t[612] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[613] = (x[11]);
  assign t[614] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[615] = (x[14]);
  assign t[616] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[617] = (x[17]);
  assign t[618] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[619] = (x[20]);
  assign t[61] = ~(t[99] | t[100]);
  assign t[620] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[621] = (x[24]);
  assign t[622] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[623] = (x[30]);
  assign t[624] = (x[25]);
  assign t[625] = (x[26]);
  assign t[626] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[627] = (x[38]);
  assign t[628] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[629] = (x[46]);
  assign t[62] = ~(t[101] ^ t[102]);
  assign t[630] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[631] = (x[52]);
  assign t[632] = (x[31]);
  assign t[633] = (x[32]);
  assign t[634] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[635] = (x[60]);
  assign t[636] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[637] = (x[68]);
  assign t[638] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[639] = (x[74]);
  assign t[63] = ~(t[103] | t[104]);
  assign t[640] = (x[23]);
  assign t[641] = (x[39]);
  assign t[642] = (x[40]);
  assign t[643] = (x[47]);
  assign t[644] = (x[48]);
  assign t[645] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[646] = (x[85]);
  assign t[647] = (x[53]);
  assign t[648] = (x[54]);
  assign t[649] = (x[29]);
  assign t[64] = ~(t[414] | t[105]);
  assign t[650] = (x[61]);
  assign t[651] = (x[62]);
  assign t[652] = (x[69]);
  assign t[653] = (x[70]);
  assign t[654] = (x[101] & ~x[102] & ~x[103] & ~x[104]) | (~x[101] & x[102] & ~x[103] & ~x[104]) | (~x[101] & ~x[102] & x[103] & ~x[104]) | (~x[101] & ~x[102] & ~x[103] & x[104]) | (x[101] & x[102] & x[103] & ~x[104]) | (x[101] & x[102] & ~x[103] & x[104]) | (x[101] & ~x[102] & x[103] & x[104]) | (~x[101] & x[102] & x[103] & x[104]);
  assign t[655] = (x[102]);
  assign t[656] = (x[75]);
  assign t[657] = (x[76]);
  assign t[658] = (x[37]);
  assign t[659] = (x[45]);
  assign t[65] = ~(t[106] ^ t[107]);
  assign t[660] = (x[86]);
  assign t[661] = (x[87]);
  assign t[662] = (x[51]);
  assign t[663] = (x[59]);
  assign t[664] = (x[67]);
  assign t[665] = (x[103]);
  assign t[666] = (x[104]);
  assign t[667] = (x[73]);
  assign t[668] = (x[84]);
  assign t[669] = (x[101]);
  assign t[66] = ~(t[415]);
  assign t[670] = (x[1]);
  assign t[671] = (x[2]);
  assign t[672] = (x[3]);
  assign t[67] = ~(t[416]);
  assign t[68] = ~(t[108] | t[109]);
  assign t[69] = ~(t[110] | t[111]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[417] | t[112]);
  assign t[71] = t[406] ? x[66] : x[65];
  assign t[72] = ~(t[30] & t[113]);
  assign t[73] = ~(t[114] | t[115]);
  assign t[74] = ~(t[418] | t[116]);
  assign t[75] = ~(t[117] | t[118]);
  assign t[76] = ~(t[119] ^ t[120]);
  assign t[77] = ~(t[121] | t[122]);
  assign t[78] = ~(t[419] | t[123]);
  assign t[79] = ~(t[124] ^ t[125]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[84]);
  assign t[81] = t[404] ? t[127] : t[126];
  assign t[82] = ~(t[128] | t[129]);
  assign t[83] = ~(t[130] & t[131]);
  assign t[84] = ~(t[406]);
  assign t[85] = t[404] ? t[133] : t[132];
  assign t[86] = ~(t[80] | t[134]);
  assign t[87] = ~(t[135]);
  assign t[88] = ~(t[420]);
  assign t[89] = ~(t[410] | t[411]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[421]);
  assign t[91] = ~(t[422]);
  assign t[92] = ~(t[136] | t[137]);
  assign t[93] = ~(t[138]);
  assign t[94] = ~(t[128]);
  assign t[95] = ~(t[139] | t[140]);
  assign t[96] = ~(t[423]);
  assign t[97] = ~(t[424]);
  assign t[98] = ~(t[141] | t[142]);
  assign t[99] = ~(t[143] | t[144]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[205] & ~t[275] & ~t[354]) | (~t[0] & t[205] & ~t[275] & ~t[354]) | (~t[0] & ~t[205] & t[275] & ~t[354]) | (~t[0] & ~t[205] & ~t[275] & t[354]) | (t[0] & t[205] & t[275] & ~t[354]) | (t[0] & t[205] & ~t[275] & t[354]) | (t[0] & ~t[205] & t[275] & t[354]) | (~t[0] & t[205] & t[275] & t[354]);
endmodule

module R2ind116(x, y);
 input [124:0] x;
 output y;

 wire [361:0] t;
  assign t[0] = t[1] ? t[2] : t[107];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[106] | t[101]);
  assign t[104] = ~(t[149]);
  assign t[105] = ~(t[150]);
  assign t[106] = ~(t[151]);
  assign t[107] = (t[152]);
  assign t[108] = (t[153]);
  assign t[109] = (t[154]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[22] : x[21];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = t[197] ^ x[5];
  assign t[153] = t[198] ^ x[11];
  assign t[154] = t[199] ^ x[14];
  assign t[155] = t[200] ^ x[17];
  assign t[156] = t[201] ^ x[20];
  assign t[157] = t[202] ^ x[28];
  assign t[158] = t[203] ^ x[36];
  assign t[159] = t[204] ^ x[39];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[205] ^ x[40];
  assign t[161] = t[206] ^ x[46];
  assign t[162] = t[207] ^ x[52];
  assign t[163] = t[208] ^ x[60];
  assign t[164] = t[209] ^ x[63];
  assign t[165] = t[210] ^ x[64];
  assign t[166] = t[211] ^ x[70];
  assign t[167] = t[212] ^ x[76];
  assign t[168] = t[213] ^ x[84];
  assign t[169] = t[214] ^ x[87];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[88];
  assign t[171] = t[216] ^ x[89];
  assign t[172] = t[217] ^ x[90];
  assign t[173] = t[218] ^ x[91];
  assign t[174] = t[219] ^ x[92];
  assign t[175] = t[220] ^ x[93];
  assign t[176] = t[221] ^ x[99];
  assign t[177] = t[222] ^ x[100];
  assign t[178] = t[223] ^ x[101];
  assign t[179] = t[224] ^ x[102];
  assign t[17] = x[7] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[103];
  assign t[181] = t[226] ^ x[104];
  assign t[182] = t[227] ^ x[110];
  assign t[183] = t[228] ^ x[111];
  assign t[184] = t[229] ^ x[112];
  assign t[185] = t[230] ^ x[113];
  assign t[186] = t[231] ^ x[114];
  assign t[187] = t[232] ^ x[115];
  assign t[188] = t[233] ^ x[116];
  assign t[189] = t[234] ^ x[117];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[118];
  assign t[191] = t[236] ^ x[119];
  assign t[192] = t[237] ^ x[120];
  assign t[193] = t[238] ^ x[121];
  assign t[194] = t[239] ^ x[122];
  assign t[195] = t[240] ^ x[123];
  assign t[196] = t[241] ^ x[124];
  assign t[197] = (~t[242] & t[243]);
  assign t[198] = (~t[244] & t[245]);
  assign t[199] = (~t[246] & t[247]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (~t[248] & t[249]);
  assign t[201] = (~t[250] & t[251]);
  assign t[202] = (~t[252] & t[253]);
  assign t[203] = (~t[254] & t[255]);
  assign t[204] = (~t[252] & t[256]);
  assign t[205] = (~t[252] & t[257]);
  assign t[206] = (~t[258] & t[259]);
  assign t[207] = (~t[260] & t[261]);
  assign t[208] = (~t[262] & t[263]);
  assign t[209] = (~t[254] & t[264]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (~t[254] & t[265]);
  assign t[211] = (~t[266] & t[267]);
  assign t[212] = (~t[268] & t[269]);
  assign t[213] = (~t[270] & t[271]);
  assign t[214] = (~t[252] & t[272]);
  assign t[215] = (~t[258] & t[273]);
  assign t[216] = (~t[258] & t[274]);
  assign t[217] = (~t[260] & t[275]);
  assign t[218] = (~t[260] & t[276]);
  assign t[219] = (~t[262] & t[277]);
  assign t[21] = x[7] ? t[33] : t[32];
  assign t[220] = (~t[262] & t[278]);
  assign t[221] = (~t[279] & t[280]);
  assign t[222] = (~t[254] & t[281]);
  assign t[223] = (~t[266] & t[282]);
  assign t[224] = (~t[266] & t[283]);
  assign t[225] = (~t[268] & t[284]);
  assign t[226] = (~t[268] & t[285]);
  assign t[227] = (~t[286] & t[287]);
  assign t[228] = (~t[270] & t[288]);
  assign t[229] = (~t[270] & t[289]);
  assign t[22] = x[7] ? t[35] : t[34];
  assign t[230] = (~t[258] & t[290]);
  assign t[231] = (~t[260] & t[291]);
  assign t[232] = (~t[262] & t[292]);
  assign t[233] = (~t[279] & t[293]);
  assign t[234] = (~t[279] & t[294]);
  assign t[235] = (~t[266] & t[295]);
  assign t[236] = (~t[268] & t[296]);
  assign t[237] = (~t[286] & t[297]);
  assign t[238] = (~t[286] & t[298]);
  assign t[239] = (~t[270] & t[299]);
  assign t[23] = ~(t[110]);
  assign t[240] = (~t[279] & t[300]);
  assign t[241] = (~t[286] & t[301]);
  assign t[242] = t[302] ^ x[4];
  assign t[243] = t[303] ^ x[5];
  assign t[244] = t[304] ^ x[10];
  assign t[245] = t[305] ^ x[11];
  assign t[246] = t[306] ^ x[13];
  assign t[247] = t[307] ^ x[14];
  assign t[248] = t[308] ^ x[16];
  assign t[249] = t[309] ^ x[17];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[310] ^ x[19];
  assign t[251] = t[311] ^ x[20];
  assign t[252] = t[312] ^ x[27];
  assign t[253] = t[313] ^ x[28];
  assign t[254] = t[314] ^ x[35];
  assign t[255] = t[315] ^ x[36];
  assign t[256] = t[316] ^ x[39];
  assign t[257] = t[317] ^ x[40];
  assign t[258] = t[318] ^ x[45];
  assign t[259] = t[319] ^ x[46];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[320] ^ x[51];
  assign t[261] = t[321] ^ x[52];
  assign t[262] = t[322] ^ x[59];
  assign t[263] = t[323] ^ x[60];
  assign t[264] = t[324] ^ x[63];
  assign t[265] = t[325] ^ x[64];
  assign t[266] = t[326] ^ x[69];
  assign t[267] = t[327] ^ x[70];
  assign t[268] = t[328] ^ x[75];
  assign t[269] = t[329] ^ x[76];
  assign t[26] = x[7] ? t[41] : t[40];
  assign t[270] = t[330] ^ x[83];
  assign t[271] = t[331] ^ x[84];
  assign t[272] = t[332] ^ x[87];
  assign t[273] = t[333] ^ x[88];
  assign t[274] = t[334] ^ x[89];
  assign t[275] = t[335] ^ x[90];
  assign t[276] = t[336] ^ x[91];
  assign t[277] = t[337] ^ x[92];
  assign t[278] = t[338] ^ x[93];
  assign t[279] = t[339] ^ x[98];
  assign t[27] = x[7] ? t[43] : t[42];
  assign t[280] = t[340] ^ x[99];
  assign t[281] = t[341] ^ x[100];
  assign t[282] = t[342] ^ x[101];
  assign t[283] = t[343] ^ x[102];
  assign t[284] = t[344] ^ x[103];
  assign t[285] = t[345] ^ x[104];
  assign t[286] = t[346] ^ x[109];
  assign t[287] = t[347] ^ x[110];
  assign t[288] = t[348] ^ x[111];
  assign t[289] = t[349] ^ x[112];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[350] ^ x[113];
  assign t[291] = t[351] ^ x[114];
  assign t[292] = t[352] ^ x[115];
  assign t[293] = t[353] ^ x[116];
  assign t[294] = t[354] ^ x[117];
  assign t[295] = t[355] ^ x[118];
  assign t[296] = t[356] ^ x[119];
  assign t[297] = t[357] ^ x[120];
  assign t[298] = t[358] ^ x[121];
  assign t[299] = t[359] ^ x[122];
  assign t[29] = t[46] | t[112];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = t[360] ^ x[123];
  assign t[301] = t[361] ^ x[124];
  assign t[302] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[303] = (x[3]);
  assign t[304] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[305] = (x[9]);
  assign t[306] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[307] = (x[12]);
  assign t[308] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[309] = (x[15]);
  assign t[30] = t[16] ? x[30] : x[29];
  assign t[310] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[311] = (x[18]);
  assign t[312] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[313] = (x[24]);
  assign t[314] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[315] = (x[32]);
  assign t[316] = (x[26]);
  assign t[317] = (x[23]);
  assign t[318] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[319] = (x[42]);
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[321] = (x[48]);
  assign t[322] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[323] = (x[56]);
  assign t[324] = (x[34]);
  assign t[325] = (x[31]);
  assign t[326] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[327] = (x[66]);
  assign t[328] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[329] = (x[72]);
  assign t[32] = ~(t[49] & t[50]);
  assign t[330] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[331] = (x[80]);
  assign t[332] = (x[25]);
  assign t[333] = (x[44]);
  assign t[334] = (x[41]);
  assign t[335] = (x[50]);
  assign t[336] = (x[47]);
  assign t[337] = (x[58]);
  assign t[338] = (x[55]);
  assign t[339] = (x[94] & ~x[95] & ~x[96] & ~x[97]) | (~x[94] & x[95] & ~x[96] & ~x[97]) | (~x[94] & ~x[95] & x[96] & ~x[97]) | (~x[94] & ~x[95] & ~x[96] & x[97]) | (x[94] & x[95] & x[96] & ~x[97]) | (x[94] & x[95] & ~x[96] & x[97]) | (x[94] & ~x[95] & x[96] & x[97]) | (~x[94] & x[95] & x[96] & x[97]);
  assign t[33] = t[51] ^ t[40];
  assign t[340] = (x[95]);
  assign t[341] = (x[33]);
  assign t[342] = (x[68]);
  assign t[343] = (x[65]);
  assign t[344] = (x[74]);
  assign t[345] = (x[71]);
  assign t[346] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[347] = (x[106]);
  assign t[348] = (x[82]);
  assign t[349] = (x[79]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[43]);
  assign t[351] = (x[49]);
  assign t[352] = (x[57]);
  assign t[353] = (x[97]);
  assign t[354] = (x[94]);
  assign t[355] = (x[67]);
  assign t[356] = (x[73]);
  assign t[357] = (x[108]);
  assign t[358] = (x[105]);
  assign t[359] = (x[81]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[96]);
  assign t[361] = (x[107]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[37] = t[58] | t[113];
  assign t[38] = t[110] ? x[38] : x[37];
  assign t[39] = ~(t[59] & t[60]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[61] & t[62]);
  assign t[41] = t[63] ^ t[64];
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[114]);
  assign t[45] = ~(t[115]);
  assign t[46] = ~(t[68] | t[44]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = t[71] | t[116];
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = ~(x[6]);
  assign t[50] = t[74] | t[117];
  assign t[51] = t[75] ? x[54] : x[53];
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = t[78] | t[118];
  assign t[54] = t[75] ? x[62] : x[61];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[119]);
  assign t[57] = ~(t[120]);
  assign t[58] = ~(t[81] | t[56]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[84] | t[121];
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = t[87] | t[122];
  assign t[63] = t[110] ? x[78] : x[77];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = t[92] | t[123];
  assign t[67] = t[110] ? x[86] : x[85];
  assign t[68] = ~(t[124]);
  assign t[69] = ~(t[125]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[126]);
  assign t[71] = ~(t[93] | t[69]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[128]);
  assign t[74] = ~(t[94] | t[72]);
  assign t[75] = ~(t[23]);
  assign t[76] = ~(t[129]);
  assign t[77] = ~(t[130]);
  assign t[78] = ~(t[95] | t[76]);
  assign t[79] = ~(t[96] & t[97]);
  assign t[7] = ~(t[108] & t[109]);
  assign t[80] = t[98] | t[131];
  assign t[81] = ~(t[132]);
  assign t[82] = ~(t[133]);
  assign t[83] = ~(t[134]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[135]);
  assign t[86] = ~(t[136]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[101] & t[102]);
  assign t[89] = t[103] | t[137];
  assign t[8] = ~(t[110] & t[111]);
  assign t[90] = ~(t[138]);
  assign t[91] = ~(t[139]);
  assign t[92] = ~(t[104] | t[90]);
  assign t[93] = ~(t[140]);
  assign t[94] = ~(t[141]);
  assign t[95] = ~(t[142]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[105] | t[96]);
  assign t[99] = ~(t[145]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [124:0] x;
 output y;

 wire [371:0] t;
  assign t[0] = t[1] ? t[2] : t[117];
  assign t[100] = ~(t[152]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[113] & t[114]);
  assign t[104] = ~(t[144] & t[143]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[156]);
  assign t[108] = ~(t[157]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[115] & t[116]);
  assign t[111] = ~(t[149] & t[148]);
  assign t[112] = ~(t[159]);
  assign t[113] = ~(t[154] & t[153]);
  assign t[114] = ~(t[160]);
  assign t[115] = ~(t[158] & t[157]);
  assign t[116] = ~(t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[21] : x[22];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = t[207] ^ x[5];
  assign t[163] = t[208] ^ x[11];
  assign t[164] = t[209] ^ x[14];
  assign t[165] = t[210] ^ x[17];
  assign t[166] = t[211] ^ x[20];
  assign t[167] = t[212] ^ x[28];
  assign t[168] = t[213] ^ x[36];
  assign t[169] = t[214] ^ x[39];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[40];
  assign t[171] = t[216] ^ x[46];
  assign t[172] = t[217] ^ x[52];
  assign t[173] = t[218] ^ x[60];
  assign t[174] = t[219] ^ x[63];
  assign t[175] = t[220] ^ x[64];
  assign t[176] = t[221] ^ x[70];
  assign t[177] = t[222] ^ x[76];
  assign t[178] = t[223] ^ x[84];
  assign t[179] = t[224] ^ x[87];
  assign t[17] = x[7] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[88];
  assign t[181] = t[226] ^ x[89];
  assign t[182] = t[227] ^ x[90];
  assign t[183] = t[228] ^ x[91];
  assign t[184] = t[229] ^ x[92];
  assign t[185] = t[230] ^ x[93];
  assign t[186] = t[231] ^ x[99];
  assign t[187] = t[232] ^ x[100];
  assign t[188] = t[233] ^ x[101];
  assign t[189] = t[234] ^ x[102];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[103];
  assign t[191] = t[236] ^ x[104];
  assign t[192] = t[237] ^ x[110];
  assign t[193] = t[238] ^ x[111];
  assign t[194] = t[239] ^ x[112];
  assign t[195] = t[240] ^ x[113];
  assign t[196] = t[241] ^ x[114];
  assign t[197] = t[242] ^ x[115];
  assign t[198] = t[243] ^ x[116];
  assign t[199] = t[244] ^ x[117];
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[245] ^ x[118];
  assign t[201] = t[246] ^ x[119];
  assign t[202] = t[247] ^ x[120];
  assign t[203] = t[248] ^ x[121];
  assign t[204] = t[249] ^ x[122];
  assign t[205] = t[250] ^ x[123];
  assign t[206] = t[251] ^ x[124];
  assign t[207] = (~t[252] & t[253]);
  assign t[208] = (~t[254] & t[255]);
  assign t[209] = (~t[256] & t[257]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (~t[258] & t[259]);
  assign t[211] = (~t[260] & t[261]);
  assign t[212] = (~t[262] & t[263]);
  assign t[213] = (~t[264] & t[265]);
  assign t[214] = (~t[262] & t[266]);
  assign t[215] = (~t[262] & t[267]);
  assign t[216] = (~t[268] & t[269]);
  assign t[217] = (~t[270] & t[271]);
  assign t[218] = (~t[272] & t[273]);
  assign t[219] = (~t[264] & t[274]);
  assign t[21] = x[7] ? t[33] : t[32];
  assign t[220] = (~t[264] & t[275]);
  assign t[221] = (~t[276] & t[277]);
  assign t[222] = (~t[278] & t[279]);
  assign t[223] = (~t[280] & t[281]);
  assign t[224] = (~t[262] & t[282]);
  assign t[225] = (~t[268] & t[283]);
  assign t[226] = (~t[268] & t[284]);
  assign t[227] = (~t[270] & t[285]);
  assign t[228] = (~t[270] & t[286]);
  assign t[229] = (~t[272] & t[287]);
  assign t[22] = x[7] ? t[35] : t[34];
  assign t[230] = (~t[272] & t[288]);
  assign t[231] = (~t[289] & t[290]);
  assign t[232] = (~t[264] & t[291]);
  assign t[233] = (~t[276] & t[292]);
  assign t[234] = (~t[276] & t[293]);
  assign t[235] = (~t[278] & t[294]);
  assign t[236] = (~t[278] & t[295]);
  assign t[237] = (~t[296] & t[297]);
  assign t[238] = (~t[280] & t[298]);
  assign t[239] = (~t[280] & t[299]);
  assign t[23] = ~(t[120]);
  assign t[240] = (~t[268] & t[300]);
  assign t[241] = (~t[270] & t[301]);
  assign t[242] = (~t[272] & t[302]);
  assign t[243] = (~t[289] & t[303]);
  assign t[244] = (~t[289] & t[304]);
  assign t[245] = (~t[276] & t[305]);
  assign t[246] = (~t[278] & t[306]);
  assign t[247] = (~t[296] & t[307]);
  assign t[248] = (~t[296] & t[308]);
  assign t[249] = (~t[280] & t[309]);
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = (~t[289] & t[310]);
  assign t[251] = (~t[296] & t[311]);
  assign t[252] = t[312] ^ x[4];
  assign t[253] = t[313] ^ x[5];
  assign t[254] = t[314] ^ x[10];
  assign t[255] = t[315] ^ x[11];
  assign t[256] = t[316] ^ x[13];
  assign t[257] = t[317] ^ x[14];
  assign t[258] = t[318] ^ x[16];
  assign t[259] = t[319] ^ x[17];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[320] ^ x[19];
  assign t[261] = t[321] ^ x[20];
  assign t[262] = t[322] ^ x[27];
  assign t[263] = t[323] ^ x[28];
  assign t[264] = t[324] ^ x[35];
  assign t[265] = t[325] ^ x[36];
  assign t[266] = t[326] ^ x[39];
  assign t[267] = t[327] ^ x[40];
  assign t[268] = t[328] ^ x[45];
  assign t[269] = t[329] ^ x[46];
  assign t[26] = x[7] ? t[41] : t[40];
  assign t[270] = t[330] ^ x[51];
  assign t[271] = t[331] ^ x[52];
  assign t[272] = t[332] ^ x[59];
  assign t[273] = t[333] ^ x[60];
  assign t[274] = t[334] ^ x[63];
  assign t[275] = t[335] ^ x[64];
  assign t[276] = t[336] ^ x[69];
  assign t[277] = t[337] ^ x[70];
  assign t[278] = t[338] ^ x[75];
  assign t[279] = t[339] ^ x[76];
  assign t[27] = x[7] ? t[43] : t[42];
  assign t[280] = t[340] ^ x[83];
  assign t[281] = t[341] ^ x[84];
  assign t[282] = t[342] ^ x[87];
  assign t[283] = t[343] ^ x[88];
  assign t[284] = t[344] ^ x[89];
  assign t[285] = t[345] ^ x[90];
  assign t[286] = t[346] ^ x[91];
  assign t[287] = t[347] ^ x[92];
  assign t[288] = t[348] ^ x[93];
  assign t[289] = t[349] ^ x[98];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[350] ^ x[99];
  assign t[291] = t[351] ^ x[100];
  assign t[292] = t[352] ^ x[101];
  assign t[293] = t[353] ^ x[102];
  assign t[294] = t[354] ^ x[103];
  assign t[295] = t[355] ^ x[104];
  assign t[296] = t[356] ^ x[109];
  assign t[297] = t[357] ^ x[110];
  assign t[298] = t[358] ^ x[111];
  assign t[299] = t[359] ^ x[112];
  assign t[29] = ~(t[46] & t[122]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = t[360] ^ x[113];
  assign t[301] = t[361] ^ x[114];
  assign t[302] = t[362] ^ x[115];
  assign t[303] = t[363] ^ x[116];
  assign t[304] = t[364] ^ x[117];
  assign t[305] = t[365] ^ x[118];
  assign t[306] = t[366] ^ x[119];
  assign t[307] = t[367] ^ x[120];
  assign t[308] = t[368] ^ x[121];
  assign t[309] = t[369] ^ x[122];
  assign t[30] = t[47] ? x[30] : x[29];
  assign t[310] = t[370] ^ x[123];
  assign t[311] = t[371] ^ x[124];
  assign t[312] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[313] = (x[2]);
  assign t[314] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[315] = (x[9]);
  assign t[316] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[317] = (x[12]);
  assign t[318] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[319] = (x[15]);
  assign t[31] = ~(t[48] & t[49]);
  assign t[320] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[321] = (x[18]);
  assign t[322] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[323] = (x[24]);
  assign t[324] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[325] = (x[32]);
  assign t[326] = (x[26]);
  assign t[327] = (x[23]);
  assign t[328] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[329] = (x[42]);
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[331] = (x[48]);
  assign t[332] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[333] = (x[56]);
  assign t[334] = (x[34]);
  assign t[335] = (x[31]);
  assign t[336] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[337] = (x[66]);
  assign t[338] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[339] = (x[72]);
  assign t[33] = t[52] ^ t[40];
  assign t[340] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[341] = (x[80]);
  assign t[342] = (x[25]);
  assign t[343] = (x[44]);
  assign t[344] = (x[41]);
  assign t[345] = (x[50]);
  assign t[346] = (x[47]);
  assign t[347] = (x[58]);
  assign t[348] = (x[55]);
  assign t[349] = (x[94] & ~x[95] & ~x[96] & ~x[97]) | (~x[94] & x[95] & ~x[96] & ~x[97]) | (~x[94] & ~x[95] & x[96] & ~x[97]) | (~x[94] & ~x[95] & ~x[96] & x[97]) | (x[94] & x[95] & x[96] & ~x[97]) | (x[94] & x[95] & ~x[96] & x[97]) | (x[94] & ~x[95] & x[96] & x[97]) | (~x[94] & x[95] & x[96] & x[97]);
  assign t[34] = ~(t[53] & t[54]);
  assign t[350] = (x[95]);
  assign t[351] = (x[33]);
  assign t[352] = (x[68]);
  assign t[353] = (x[65]);
  assign t[354] = (x[74]);
  assign t[355] = (x[71]);
  assign t[356] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[357] = (x[106]);
  assign t[358] = (x[82]);
  assign t[359] = (x[79]);
  assign t[35] = t[55] ^ t[56];
  assign t[360] = (x[43]);
  assign t[361] = (x[49]);
  assign t[362] = (x[57]);
  assign t[363] = (x[97]);
  assign t[364] = (x[94]);
  assign t[365] = (x[67]);
  assign t[366] = (x[73]);
  assign t[367] = (x[108]);
  assign t[368] = (x[105]);
  assign t[369] = (x[81]);
  assign t[36] = ~(t[57] & t[58]);
  assign t[370] = (x[96]);
  assign t[371] = (x[107]);
  assign t[37] = ~(t[59] & t[123]);
  assign t[38] = t[120] ? x[38] : x[37];
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[62] & t[63]);
  assign t[41] = t[64] ^ t[65];
  assign t[42] = ~(t[66] & t[67]);
  assign t[43] = t[68] ^ t[42];
  assign t[44] = ~(t[124]);
  assign t[45] = ~(t[125]);
  assign t[46] = ~(t[69] & t[70]);
  assign t[47] = ~(t[23]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[73] & t[126]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = ~(t[76] & t[127]);
  assign t[52] = t[16] ? x[54] : x[53];
  assign t[53] = ~(t[77] & t[78]);
  assign t[54] = ~(t[79] & t[128]);
  assign t[55] = t[16] ? x[62] : x[61];
  assign t[56] = ~(t[80] & t[81]);
  assign t[57] = ~(t[129]);
  assign t[58] = ~(t[130]);
  assign t[59] = ~(t[82] & t[83]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = ~(t[86] & t[131]);
  assign t[62] = ~(t[87] & t[88]);
  assign t[63] = ~(t[89] & t[132]);
  assign t[64] = t[120] ? x[78] : x[77];
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = ~(t[92] & t[93]);
  assign t[67] = ~(t[94] & t[133]);
  assign t[68] = t[120] ? x[86] : x[85];
  assign t[69] = ~(t[125] & t[124]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[134]);
  assign t[71] = ~(t[135]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[95] & t[96]);
  assign t[74] = ~(t[137]);
  assign t[75] = ~(t[138]);
  assign t[76] = ~(t[97] & t[98]);
  assign t[77] = ~(t[139]);
  assign t[78] = ~(t[140]);
  assign t[79] = ~(t[99] & t[100]);
  assign t[7] = ~(t[118] & t[119]);
  assign t[80] = ~(t[101] & t[102]);
  assign t[81] = ~(t[103] & t[141]);
  assign t[82] = ~(t[130] & t[129]);
  assign t[83] = ~(t[142]);
  assign t[84] = ~(t[143]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[104] & t[105]);
  assign t[87] = ~(t[145]);
  assign t[88] = ~(t[146]);
  assign t[89] = ~(t[106] & t[107]);
  assign t[8] = ~(t[120] & t[121]);
  assign t[90] = ~(t[108] & t[109]);
  assign t[91] = ~(t[110] & t[147]);
  assign t[92] = ~(t[148]);
  assign t[93] = ~(t[149]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[136] & t[135]);
  assign t[96] = ~(t[150]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[151]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [114:0] x;
 output y;

 wire [302:0] t;
  assign t[0] = t[1] ? t[2] : t[98];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[16] ? x[21] : x[22];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = t[168] ^ x[5];
  assign t[134] = t[169] ^ x[11];
  assign t[135] = t[170] ^ x[14];
  assign t[136] = t[171] ^ x[17];
  assign t[137] = t[172] ^ x[20];
  assign t[138] = t[173] ^ x[28];
  assign t[139] = t[174] ^ x[29];
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = t[175] ^ x[37];
  assign t[141] = t[176] ^ x[38];
  assign t[142] = t[177] ^ x[41];
  assign t[143] = t[178] ^ x[47];
  assign t[144] = t[179] ^ x[48];
  assign t[145] = t[180] ^ x[54];
  assign t[146] = t[181] ^ x[55];
  assign t[147] = t[182] ^ x[63];
  assign t[148] = t[183] ^ x[64];
  assign t[149] = t[184] ^ x[67];
  assign t[14] = x[7] ? t[20] : t[19];
  assign t[150] = t[185] ^ x[73];
  assign t[151] = t[186] ^ x[74];
  assign t[152] = t[187] ^ x[80];
  assign t[153] = t[188] ^ x[81];
  assign t[154] = t[189] ^ x[89];
  assign t[155] = t[190] ^ x[90];
  assign t[156] = t[191] ^ x[93];
  assign t[157] = t[192] ^ x[94];
  assign t[158] = t[193] ^ x[95];
  assign t[159] = t[194] ^ x[101];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[195] ^ x[102];
  assign t[161] = t[196] ^ x[103];
  assign t[162] = t[197] ^ x[104];
  assign t[163] = t[198] ^ x[105];
  assign t[164] = t[199] ^ x[111];
  assign t[165] = t[200] ^ x[112];
  assign t[166] = t[201] ^ x[113];
  assign t[167] = t[202] ^ x[114];
  assign t[168] = (~t[203] & t[204]);
  assign t[169] = (~t[205] & t[206]);
  assign t[16] = ~(t[23]);
  assign t[170] = (~t[207] & t[208]);
  assign t[171] = (~t[209] & t[210]);
  assign t[172] = (~t[211] & t[212]);
  assign t[173] = (~t[213] & t[214]);
  assign t[174] = (~t[213] & t[215]);
  assign t[175] = (~t[216] & t[217]);
  assign t[176] = (~t[216] & t[218]);
  assign t[177] = (~t[213] & t[219]);
  assign t[178] = (~t[220] & t[221]);
  assign t[179] = (~t[220] & t[222]);
  assign t[17] = x[7] ? t[25] : t[24];
  assign t[180] = (~t[223] & t[224]);
  assign t[181] = (~t[223] & t[225]);
  assign t[182] = (~t[226] & t[227]);
  assign t[183] = (~t[226] & t[228]);
  assign t[184] = (~t[216] & t[229]);
  assign t[185] = (~t[230] & t[231]);
  assign t[186] = (~t[230] & t[232]);
  assign t[187] = (~t[233] & t[234]);
  assign t[188] = (~t[233] & t[235]);
  assign t[189] = (~t[236] & t[237]);
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = (~t[236] & t[238]);
  assign t[191] = (~t[220] & t[239]);
  assign t[192] = (~t[223] & t[240]);
  assign t[193] = (~t[226] & t[241]);
  assign t[194] = (~t[242] & t[243]);
  assign t[195] = (~t[242] & t[244]);
  assign t[196] = (~t[230] & t[245]);
  assign t[197] = (~t[233] & t[246]);
  assign t[198] = (~t[236] & t[247]);
  assign t[199] = (~t[248] & t[249]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (~t[248] & t[250]);
  assign t[201] = (~t[242] & t[251]);
  assign t[202] = (~t[248] & t[252]);
  assign t[203] = t[253] ^ x[4];
  assign t[204] = t[254] ^ x[5];
  assign t[205] = t[255] ^ x[10];
  assign t[206] = t[256] ^ x[11];
  assign t[207] = t[257] ^ x[13];
  assign t[208] = t[258] ^ x[14];
  assign t[209] = t[259] ^ x[16];
  assign t[20] = t[30] ^ t[31];
  assign t[210] = t[260] ^ x[17];
  assign t[211] = t[261] ^ x[19];
  assign t[212] = t[262] ^ x[20];
  assign t[213] = t[263] ^ x[27];
  assign t[214] = t[264] ^ x[28];
  assign t[215] = t[265] ^ x[29];
  assign t[216] = t[266] ^ x[36];
  assign t[217] = t[267] ^ x[37];
  assign t[218] = t[268] ^ x[38];
  assign t[219] = t[269] ^ x[41];
  assign t[21] = x[7] ? t[33] : t[32];
  assign t[220] = t[270] ^ x[46];
  assign t[221] = t[271] ^ x[47];
  assign t[222] = t[272] ^ x[48];
  assign t[223] = t[273] ^ x[53];
  assign t[224] = t[274] ^ x[54];
  assign t[225] = t[275] ^ x[55];
  assign t[226] = t[276] ^ x[62];
  assign t[227] = t[277] ^ x[63];
  assign t[228] = t[278] ^ x[64];
  assign t[229] = t[279] ^ x[67];
  assign t[22] = x[7] ? t[35] : t[34];
  assign t[230] = t[280] ^ x[72];
  assign t[231] = t[281] ^ x[73];
  assign t[232] = t[282] ^ x[74];
  assign t[233] = t[283] ^ x[79];
  assign t[234] = t[284] ^ x[80];
  assign t[235] = t[285] ^ x[81];
  assign t[236] = t[286] ^ x[88];
  assign t[237] = t[287] ^ x[89];
  assign t[238] = t[288] ^ x[90];
  assign t[239] = t[289] ^ x[93];
  assign t[23] = ~(t[101]);
  assign t[240] = t[290] ^ x[94];
  assign t[241] = t[291] ^ x[95];
  assign t[242] = t[292] ^ x[100];
  assign t[243] = t[293] ^ x[101];
  assign t[244] = t[294] ^ x[102];
  assign t[245] = t[295] ^ x[103];
  assign t[246] = t[296] ^ x[104];
  assign t[247] = t[297] ^ x[105];
  assign t[248] = t[298] ^ x[110];
  assign t[249] = t[299] ^ x[111];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[300] ^ x[112];
  assign t[251] = t[301] ^ x[113];
  assign t[252] = t[302] ^ x[114];
  assign t[253] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[254] = (x[1]);
  assign t[255] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[256] = (x[9]);
  assign t[257] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[258] = (x[12]);
  assign t[259] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[25] = t[38] ^ t[39];
  assign t[260] = (x[15]);
  assign t[261] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[262] = (x[18]);
  assign t[263] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[264] = (x[25]);
  assign t[265] = (x[23]);
  assign t[266] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[267] = (x[34]);
  assign t[268] = (x[32]);
  assign t[269] = (x[26]);
  assign t[26] = x[7] ? t[41] : t[40];
  assign t[270] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[271] = (x[44]);
  assign t[272] = (x[42]);
  assign t[273] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[274] = (x[51]);
  assign t[275] = (x[49]);
  assign t[276] = (x[58] & ~x[59] & ~x[60] & ~x[61]) | (~x[58] & x[59] & ~x[60] & ~x[61]) | (~x[58] & ~x[59] & x[60] & ~x[61]) | (~x[58] & ~x[59] & ~x[60] & x[61]) | (x[58] & x[59] & x[60] & ~x[61]) | (x[58] & x[59] & ~x[60] & x[61]) | (x[58] & ~x[59] & x[60] & x[61]) | (~x[58] & x[59] & x[60] & x[61]);
  assign t[277] = (x[60]);
  assign t[278] = (x[58]);
  assign t[279] = (x[35]);
  assign t[27] = x[7] ? t[43] : t[42];
  assign t[280] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[281] = (x[70]);
  assign t[282] = (x[68]);
  assign t[283] = (x[75] & ~x[76] & ~x[77] & ~x[78]) | (~x[75] & x[76] & ~x[77] & ~x[78]) | (~x[75] & ~x[76] & x[77] & ~x[78]) | (~x[75] & ~x[76] & ~x[77] & x[78]) | (x[75] & x[76] & x[77] & ~x[78]) | (x[75] & x[76] & ~x[77] & x[78]) | (x[75] & ~x[76] & x[77] & x[78]) | (~x[75] & x[76] & x[77] & x[78]);
  assign t[284] = (x[77]);
  assign t[285] = (x[75]);
  assign t[286] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[287] = (x[86]);
  assign t[288] = (x[84]);
  assign t[289] = (x[45]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[290] = (x[52]);
  assign t[291] = (x[61]);
  assign t[292] = (x[96] & ~x[97] & ~x[98] & ~x[99]) | (~x[96] & x[97] & ~x[98] & ~x[99]) | (~x[96] & ~x[97] & x[98] & ~x[99]) | (~x[96] & ~x[97] & ~x[98] & x[99]) | (x[96] & x[97] & x[98] & ~x[99]) | (x[96] & x[97] & ~x[98] & x[99]) | (x[96] & ~x[97] & x[98] & x[99]) | (~x[96] & x[97] & x[98] & x[99]);
  assign t[293] = (x[98]);
  assign t[294] = (x[96]);
  assign t[295] = (x[71]);
  assign t[296] = (x[78]);
  assign t[297] = (x[87]);
  assign t[298] = (x[106] & ~x[107] & ~x[108] & ~x[109]) | (~x[106] & x[107] & ~x[108] & ~x[109]) | (~x[106] & ~x[107] & x[108] & ~x[109]) | (~x[106] & ~x[107] & ~x[108] & x[109]) | (x[106] & x[107] & x[108] & ~x[109]) | (x[106] & x[107] & ~x[108] & x[109]) | (x[106] & ~x[107] & x[108] & x[109]) | (~x[106] & x[107] & x[108] & x[109]);
  assign t[299] = (x[108]);
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = (x[106]);
  assign t[301] = (x[99]);
  assign t[302] = (x[109]);
  assign t[30] = t[46] ? x[31] : x[30];
  assign t[31] = ~(t[47] & t[48]);
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = t[51] ^ t[42];
  assign t[34] = ~(t[52] & t[53]);
  assign t[35] = t[54] ^ t[55];
  assign t[36] = ~(t[105] & t[56]);
  assign t[37] = ~(t[106] & t[57]);
  assign t[38] = t[101] ? x[40] : x[39];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[40];
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[107]);
  assign t[45] = ~(t[107] & t[67]);
  assign t[46] = ~(t[23]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = t[72] ? x[57] : x[56];
  assign t[52] = ~(t[112] & t[73]);
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = t[72] ? x[66] : x[65];
  assign t[55] = ~(t[75] & t[76]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[114] & t[77]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = t[101] ? x[83] : x[82];
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = ~(t[120] & t[83]);
  assign t[65] = t[101] ? x[92] : x[91];
  assign t[66] = ~(t[84] & t[85]);
  assign t[67] = ~(t[103]);
  assign t[68] = ~(t[121]);
  assign t[69] = ~(t[121] & t[86]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[122]);
  assign t[71] = ~(t[122] & t[87]);
  assign t[72] = ~(t[23]);
  assign t[73] = ~(t[123]);
  assign t[74] = ~(t[123] & t[88]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[105]);
  assign t[78] = ~(t[126]);
  assign t[79] = ~(t[126] & t[91]);
  assign t[7] = ~(t[99] & t[100]);
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[131]);
  assign t[8] = ~(t[101] & t[102]);
  assign t[90] = ~(t[131] & t[96]);
  assign t[91] = ~(t[115]);
  assign t[92] = ~(t[117]);
  assign t[93] = ~(t[119]);
  assign t[94] = ~(t[132]);
  assign t[95] = ~(t[132] & t[97]);
  assign t[96] = ~(t[124]);
  assign t[97] = ~(t[129]);
  assign t[98] = (t[133]);
  assign t[99] = (t[134]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [124:0] x;
 output y;

 wire [459:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = ~(t[227] | t[145]);
  assign t[101] = t[146] ? x[91] : x[90];
  assign t[102] = ~(t[147] & t[83]);
  assign t[103] = ~(t[228]);
  assign t[104] = ~(t[229]);
  assign t[105] = ~(t[148] | t[149]);
  assign t[106] = t[146] ? x[95] : x[94];
  assign t[107] = ~(t[150] & t[151]);
  assign t[108] = ~(t[230]);
  assign t[109] = ~(t[217] | t[218]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[232]);
  assign t[112] = ~(t[152] | t[153]);
  assign t[113] = ~(t[154] | t[155]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[234]);
  assign t[116] = ~(t[156] | t[157]);
  assign t[117] = ~(t[158] | t[159]);
  assign t[118] = ~(t[235] | t[160]);
  assign t[119] = t[93] ? x[108] : x[107];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[161] & t[162]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[237]);
  assign t[123] = ~(t[163] | t[164]);
  assign t[124] = t[208] ? x[112] : x[111];
  assign t[125] = t[165] | t[166];
  assign t[126] = ~(t[167] & t[209]);
  assign t[127] = ~(t[168] & t[169]);
  assign t[128] = ~(t[80] | t[170]);
  assign t[129] = ~(t[80] | t[171]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[209] & t[172];
  assign t[131] = t[168] | t[167];
  assign t[132] = ~(x[7] & t[173]);
  assign t[133] = ~(t[174] & t[169]);
  assign t[134] = t[206] ? t[176] : t[175];
  assign t[135] = ~(t[172] & t[177]);
  assign t[136] = ~(t[238]);
  assign t[137] = ~(t[223] | t[224]);
  assign t[138] = ~(t[208]);
  assign t[139] = ~(t[113]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[80] | t[178]);
  assign t[141] = ~(t[239]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[240]);
  assign t[144] = ~(t[241]);
  assign t[145] = ~(t[179] | t[180]);
  assign t[146] = ~(t[138]);
  assign t[147] = ~(t[165] | t[181]);
  assign t[148] = ~(t[242]);
  assign t[149] = ~(t[228] | t[229]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[128] | t[182]);
  assign t[151] = ~(t[183] & t[184]);
  assign t[152] = ~(t[243]);
  assign t[153] = ~(t[231] | t[232]);
  assign t[154] = ~(t[80] | t[185]);
  assign t[155] = ~(t[80] | t[186]);
  assign t[156] = ~(t[244]);
  assign t[157] = ~(t[233] | t[234]);
  assign t[158] = ~(t[245]);
  assign t[159] = ~(t[246]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[187] | t[188]);
  assign t[161] = ~(t[165] | t[189]);
  assign t[162] = ~(t[48]);
  assign t[163] = ~(t[247]);
  assign t[164] = ~(t[236] | t[237]);
  assign t[165] = ~(t[135] & t[151]);
  assign t[166] = ~(t[190] & t[191]);
  assign t[167] = x[7] & t[207];
  assign t[168] = ~(x[7] | t[207]);
  assign t[169] = ~(t[209]);
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = t[206] ? t[126] : t[127];
  assign t[171] = t[206] ? t[132] : t[192];
  assign t[172] = ~(t[84] | t[206]);
  assign t[173] = ~(t[207] | t[209]);
  assign t[174] = ~(x[7] | t[193]);
  assign t[175] = ~(t[167] & t[169]);
  assign t[176] = ~(t[168] & t[209]);
  assign t[177] = ~(t[192] & t[194]);
  assign t[178] = t[206] ? t[192] : t[132];
  assign t[179] = ~(t[248]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[240] | t[241]);
  assign t[181] = t[140] | t[86];
  assign t[182] = ~(t[195] & t[196]);
  assign t[183] = ~(t[207] | t[169]);
  assign t[184] = t[80] & t[206];
  assign t[185] = t[206] ? t[194] : t[133];
  assign t[186] = t[206] ? t[175] : t[176];
  assign t[187] = ~(t[249]);
  assign t[188] = ~(t[245] | t[246]);
  assign t[189] = ~(t[197] & t[198]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[48] | t[86]);
  assign t[191] = ~(t[129] | t[155]);
  assign t[192] = ~(t[209] & t[174]);
  assign t[193] = ~(t[207]);
  assign t[194] = ~(x[7] & t[183]);
  assign t[195] = ~(t[199] | t[200]);
  assign t[196] = ~(t[84] & t[201]);
  assign t[197] = ~(t[50]);
  assign t[198] = t[84] | t[202];
  assign t[199] = ~(t[84] | t[203]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[80] | t[204]);
  assign t[201] = ~(t[132] & t[192]);
  assign t[202] = t[206] ? t[132] : t[133];
  assign t[203] = t[206] ? t[127] : t[175];
  assign t[204] = t[206] ? t[133] : t[194];
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[208] ? x[9] : x[10];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[32] | t[33]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[34] ^ t[35]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[295] ^ x[5];
  assign t[251] = t[296] ^ x[13];
  assign t[252] = t[297] ^ x[16];
  assign t[253] = t[298] ^ x[19];
  assign t[254] = t[299] ^ x[22];
  assign t[255] = t[300] ^ x[28];
  assign t[256] = t[301] ^ x[34];
  assign t[257] = t[302] ^ x[35];
  assign t[258] = t[303] ^ x[36];
  assign t[259] = t[304] ^ x[42];
  assign t[25] = x[7] ? t[39] : t[38];
  assign t[260] = t[305] ^ x[50];
  assign t[261] = t[306] ^ x[56];
  assign t[262] = t[307] ^ x[57];
  assign t[263] = t[308] ^ x[58];
  assign t[264] = t[309] ^ x[64];
  assign t[265] = t[310] ^ x[72];
  assign t[266] = t[311] ^ x[78];
  assign t[267] = t[312] ^ x[79];
  assign t[268] = t[313] ^ x[80];
  assign t[269] = t[314] ^ x[81];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[315] ^ x[82];
  assign t[271] = t[316] ^ x[83];
  assign t[272] = t[317] ^ x[89];
  assign t[273] = t[318] ^ x[92];
  assign t[274] = t[319] ^ x[93];
  assign t[275] = t[320] ^ x[96];
  assign t[276] = t[321] ^ x[97];
  assign t[277] = t[322] ^ x[98];
  assign t[278] = t[323] ^ x[99];
  assign t[279] = t[324] ^ x[100];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[325] ^ x[106];
  assign t[281] = t[326] ^ x[109];
  assign t[282] = t[327] ^ x[110];
  assign t[283] = t[328] ^ x[113];
  assign t[284] = t[329] ^ x[114];
  assign t[285] = t[330] ^ x[115];
  assign t[286] = t[331] ^ x[116];
  assign t[287] = t[332] ^ x[117];
  assign t[288] = t[333] ^ x[118];
  assign t[289] = t[334] ^ x[119];
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = t[335] ^ x[120];
  assign t[291] = t[336] ^ x[121];
  assign t[292] = t[337] ^ x[122];
  assign t[293] = t[338] ^ x[123];
  assign t[294] = t[339] ^ x[124];
  assign t[295] = (~t[340] & t[341]);
  assign t[296] = (~t[342] & t[343]);
  assign t[297] = (~t[344] & t[345]);
  assign t[298] = (~t[346] & t[347]);
  assign t[299] = (~t[348] & t[349]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[350] & t[351]);
  assign t[301] = (~t[352] & t[353]);
  assign t[302] = (~t[350] & t[354]);
  assign t[303] = (~t[350] & t[355]);
  assign t[304] = (~t[356] & t[357]);
  assign t[305] = (~t[358] & t[359]);
  assign t[306] = (~t[360] & t[361]);
  assign t[307] = (~t[352] & t[362]);
  assign t[308] = (~t[352] & t[363]);
  assign t[309] = (~t[364] & t[365]);
  assign t[30] = ~(t[48] | t[49]);
  assign t[310] = (~t[366] & t[367]);
  assign t[311] = (~t[368] & t[369]);
  assign t[312] = (~t[350] & t[370]);
  assign t[313] = (~t[356] & t[371]);
  assign t[314] = (~t[356] & t[372]);
  assign t[315] = (~t[358] & t[373]);
  assign t[316] = (~t[358] & t[374]);
  assign t[317] = (~t[375] & t[376]);
  assign t[318] = (~t[360] & t[377]);
  assign t[319] = (~t[360] & t[378]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (~t[352] & t[379]);
  assign t[321] = (~t[364] & t[380]);
  assign t[322] = (~t[364] & t[381]);
  assign t[323] = (~t[366] & t[382]);
  assign t[324] = (~t[366] & t[383]);
  assign t[325] = (~t[384] & t[385]);
  assign t[326] = (~t[368] & t[386]);
  assign t[327] = (~t[368] & t[387]);
  assign t[328] = (~t[356] & t[388]);
  assign t[329] = (~t[358] & t[389]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (~t[375] & t[390]);
  assign t[331] = (~t[375] & t[391]);
  assign t[332] = (~t[360] & t[392]);
  assign t[333] = (~t[364] & t[393]);
  assign t[334] = (~t[366] & t[394]);
  assign t[335] = (~t[384] & t[395]);
  assign t[336] = (~t[384] & t[396]);
  assign t[337] = (~t[368] & t[397]);
  assign t[338] = (~t[375] & t[398]);
  assign t[339] = (~t[384] & t[399]);
  assign t[33] = ~(t[210] | t[54]);
  assign t[340] = t[400] ^ x[4];
  assign t[341] = t[401] ^ x[5];
  assign t[342] = t[402] ^ x[12];
  assign t[343] = t[403] ^ x[13];
  assign t[344] = t[404] ^ x[15];
  assign t[345] = t[405] ^ x[16];
  assign t[346] = t[406] ^ x[18];
  assign t[347] = t[407] ^ x[19];
  assign t[348] = t[408] ^ x[21];
  assign t[349] = t[409] ^ x[22];
  assign t[34] = ~(t[55] | t[56]);
  assign t[350] = t[410] ^ x[27];
  assign t[351] = t[411] ^ x[28];
  assign t[352] = t[412] ^ x[33];
  assign t[353] = t[413] ^ x[34];
  assign t[354] = t[414] ^ x[35];
  assign t[355] = t[415] ^ x[36];
  assign t[356] = t[416] ^ x[41];
  assign t[357] = t[417] ^ x[42];
  assign t[358] = t[418] ^ x[49];
  assign t[359] = t[419] ^ x[50];
  assign t[35] = ~(t[57] ^ t[58]);
  assign t[360] = t[420] ^ x[55];
  assign t[361] = t[421] ^ x[56];
  assign t[362] = t[422] ^ x[57];
  assign t[363] = t[423] ^ x[58];
  assign t[364] = t[424] ^ x[63];
  assign t[365] = t[425] ^ x[64];
  assign t[366] = t[426] ^ x[71];
  assign t[367] = t[427] ^ x[72];
  assign t[368] = t[428] ^ x[77];
  assign t[369] = t[429] ^ x[78];
  assign t[36] = ~(t[59] | t[60]);
  assign t[370] = t[430] ^ x[79];
  assign t[371] = t[431] ^ x[80];
  assign t[372] = t[432] ^ x[81];
  assign t[373] = t[433] ^ x[82];
  assign t[374] = t[434] ^ x[83];
  assign t[375] = t[435] ^ x[88];
  assign t[376] = t[436] ^ x[89];
  assign t[377] = t[437] ^ x[92];
  assign t[378] = t[438] ^ x[93];
  assign t[379] = t[439] ^ x[96];
  assign t[37] = ~(t[61] ^ t[62]);
  assign t[380] = t[440] ^ x[97];
  assign t[381] = t[441] ^ x[98];
  assign t[382] = t[442] ^ x[99];
  assign t[383] = t[443] ^ x[100];
  assign t[384] = t[444] ^ x[105];
  assign t[385] = t[445] ^ x[106];
  assign t[386] = t[446] ^ x[109];
  assign t[387] = t[447] ^ x[110];
  assign t[388] = t[448] ^ x[113];
  assign t[389] = t[449] ^ x[114];
  assign t[38] = ~(t[63] | t[64]);
  assign t[390] = t[450] ^ x[115];
  assign t[391] = t[451] ^ x[116];
  assign t[392] = t[452] ^ x[117];
  assign t[393] = t[453] ^ x[118];
  assign t[394] = t[454] ^ x[119];
  assign t[395] = t[455] ^ x[120];
  assign t[396] = t[456] ^ x[121];
  assign t[397] = t[457] ^ x[122];
  assign t[398] = t[458] ^ x[123];
  assign t[399] = t[459] ^ x[124];
  assign t[39] = ~(t[44] ^ t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[401] = (x[0]);
  assign t[402] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[403] = (x[11]);
  assign t[404] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[405] = (x[14]);
  assign t[406] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[407] = (x[17]);
  assign t[408] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[409] = (x[20]);
  assign t[40] = ~(t[66] | t[67]);
  assign t[410] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[411] = (x[24]);
  assign t[412] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[413] = (x[30]);
  assign t[414] = (x[25]);
  assign t[415] = (x[26]);
  assign t[416] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[417] = (x[38]);
  assign t[418] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[419] = (x[46]);
  assign t[41] = ~(t[211] | t[68]);
  assign t[420] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[421] = (x[52]);
  assign t[422] = (x[31]);
  assign t[423] = (x[32]);
  assign t[424] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[425] = (x[60]);
  assign t[426] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[427] = (x[68]);
  assign t[428] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[429] = (x[74]);
  assign t[42] = ~(t[69] | t[70]);
  assign t[430] = (x[23]);
  assign t[431] = (x[39]);
  assign t[432] = (x[40]);
  assign t[433] = (x[47]);
  assign t[434] = (x[48]);
  assign t[435] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[436] = (x[85]);
  assign t[437] = (x[53]);
  assign t[438] = (x[54]);
  assign t[439] = (x[29]);
  assign t[43] = ~(t[71] ^ t[72]);
  assign t[440] = (x[61]);
  assign t[441] = (x[62]);
  assign t[442] = (x[69]);
  assign t[443] = (x[70]);
  assign t[444] = (x[101] & ~x[102] & ~x[103] & ~x[104]) | (~x[101] & x[102] & ~x[103] & ~x[104]) | (~x[101] & ~x[102] & x[103] & ~x[104]) | (~x[101] & ~x[102] & ~x[103] & x[104]) | (x[101] & x[102] & x[103] & ~x[104]) | (x[101] & x[102] & ~x[103] & x[104]) | (x[101] & ~x[102] & x[103] & x[104]) | (~x[101] & x[102] & x[103] & x[104]);
  assign t[445] = (x[102]);
  assign t[446] = (x[75]);
  assign t[447] = (x[76]);
  assign t[448] = (x[37]);
  assign t[449] = (x[45]);
  assign t[44] = ~(t[73] | t[74]);
  assign t[450] = (x[86]);
  assign t[451] = (x[87]);
  assign t[452] = (x[51]);
  assign t[453] = (x[59]);
  assign t[454] = (x[67]);
  assign t[455] = (x[103]);
  assign t[456] = (x[104]);
  assign t[457] = (x[73]);
  assign t[458] = (x[84]);
  assign t[459] = (x[101]);
  assign t[45] = ~(t[75] ^ t[76]);
  assign t[46] = ~(t[77] | t[78]);
  assign t[47] = ~(t[46] ^ t[79]);
  assign t[48] = ~(t[80] | t[81]);
  assign t[49] = ~(t[82] & t[83]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[84] | t[85]);
  assign t[51] = t[86] | t[87];
  assign t[52] = ~(t[212]);
  assign t[53] = ~(t[213]);
  assign t[54] = ~(t[88] | t[89]);
  assign t[55] = ~(t[90] | t[91]);
  assign t[56] = ~(t[214] | t[92]);
  assign t[57] = t[93] ? x[44] : x[43];
  assign t[58] = ~(t[94] & t[95]);
  assign t[59] = ~(t[96] | t[97]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[215] | t[98]);
  assign t[61] = ~(t[99] | t[100]);
  assign t[62] = ~(t[101] ^ t[102]);
  assign t[63] = ~(t[103] | t[104]);
  assign t[64] = ~(t[216] | t[105]);
  assign t[65] = ~(t[106] ^ t[107]);
  assign t[66] = ~(t[217]);
  assign t[67] = ~(t[218]);
  assign t[68] = ~(t[108] | t[109]);
  assign t[69] = ~(t[110] | t[111]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[219] | t[112]);
  assign t[71] = t[208] ? x[66] : x[65];
  assign t[72] = ~(t[30] & t[113]);
  assign t[73] = ~(t[114] | t[115]);
  assign t[74] = ~(t[220] | t[116]);
  assign t[75] = ~(t[117] | t[118]);
  assign t[76] = ~(t[119] ^ t[120]);
  assign t[77] = ~(t[121] | t[122]);
  assign t[78] = ~(t[221] | t[123]);
  assign t[79] = ~(t[124] ^ t[125]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[84]);
  assign t[81] = t[206] ? t[127] : t[126];
  assign t[82] = ~(t[128] | t[129]);
  assign t[83] = ~(t[130] & t[131]);
  assign t[84] = ~(t[208]);
  assign t[85] = t[206] ? t[133] : t[132];
  assign t[86] = ~(t[80] | t[134]);
  assign t[87] = ~(t[135]);
  assign t[88] = ~(t[222]);
  assign t[89] = ~(t[212] | t[213]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[223]);
  assign t[91] = ~(t[224]);
  assign t[92] = ~(t[136] | t[137]);
  assign t[93] = ~(t[138]);
  assign t[94] = ~(t[128]);
  assign t[95] = ~(t[139] | t[140]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[226]);
  assign t[98] = ~(t[141] | t[142]);
  assign t[99] = ~(t[143] | t[144]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [112:0] x;
 output y;

 wire [440:0] t;
  assign t[0] = t[1] ? t[2] : t[259];
  assign t[100] = ~(t[283]);
  assign t[101] = ~(t[276] | t[277]);
  assign t[102] = ~(t[284]);
  assign t[103] = ~(t[285]);
  assign t[104] = ~(t[119] | t[120]);
  assign t[105] = ~(t[121] | t[57]);
  assign t[106] = ~(x[7] | t[122]);
  assign t[107] = ~(t[123] & t[263]);
  assign t[108] = ~(t[124] & t[83]);
  assign t[109] = ~(t[123] & t[83]);
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = ~(t[124] & t[263]);
  assign t[111] = ~(x[7] & t[125]);
  assign t[112] = ~(t[117]);
  assign t[113] = t[80] | t[126];
  assign t[114] = ~(t[286]);
  assign t[115] = ~(t[281] | t[282]);
  assign t[116] = ~(t[127] & t[128]);
  assign t[117] = ~(t[80] | t[129]);
  assign t[118] = t[55] | t[130];
  assign t[119] = ~(t[287]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = ~(t[284] | t[285]);
  assign t[121] = ~(t[84] | t[131]);
  assign t[122] = ~(t[261]);
  assign t[123] = x[7] & t[261];
  assign t[124] = ~(x[7] | t[261]);
  assign t[125] = ~(t[261] | t[263]);
  assign t[126] = t[260] ? t[111] : t[132];
  assign t[127] = ~(t[133] | t[56]);
  assign t[128] = ~(t[134] & t[135]);
  assign t[129] = t[260] ? t[132] : t[111];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = ~(t[31]);
  assign t[131] = t[260] ? t[82] : t[132];
  assign t[132] = ~(t[106] & t[83]);
  assign t[133] = ~(t[84] | t[136]);
  assign t[134] = t[263] & t[50];
  assign t[135] = t[124] | t[123];
  assign t[136] = t[260] ? t[107] : t[108];
  assign t[137] = t[1] ? t[138] : t[288];
  assign t[138] = x[6] ? t[140] : t[139];
  assign t[139] = x[7] ? t[142] : t[141];
  assign t[13] = x[7] ? t[18] : t[17];
  assign t[140] = t[143] ^ x[84];
  assign t[141] = t[144] ^ t[142];
  assign t[142] = ~(t[145] ^ t[146]);
  assign t[143] = x[85] ^ x[86];
  assign t[144] = t[262] ? x[86] : x[85];
  assign t[145] = x[7] ? t[148] : t[147];
  assign t[146] = ~(t[149] ^ t[150]);
  assign t[147] = ~(t[151] & t[152]);
  assign t[148] = t[153] ^ t[154];
  assign t[149] = x[7] ? t[156] : t[155];
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = x[7] ? t[158] : t[157];
  assign t[151] = ~(t[265] & t[36]);
  assign t[152] = ~(t[270] & t[159]);
  assign t[153] = t[262] ? x[88] : x[87];
  assign t[154] = ~(t[160] & t[161]);
  assign t[155] = ~(t[162] & t[163]);
  assign t[156] = t[164] ^ t[165];
  assign t[157] = ~(t[166] & t[167]);
  assign t[158] = t[168] ^ t[169];
  assign t[159] = ~(t[266] & t[35]);
  assign t[15] = t[262] ? x[22] : x[21];
  assign t[160] = ~(t[271] & t[61]);
  assign t[161] = ~(t[279] & t[170]);
  assign t[162] = ~(t[276] & t[74]);
  assign t[163] = ~(t[283] & t[171]);
  assign t[164] = t[262] ? x[90] : x[89];
  assign t[165] = ~(t[172] & t[173]);
  assign t[166] = ~(t[273] & t[67]);
  assign t[167] = ~(t[280] & t[174]);
  assign t[168] = t[175] ? x[92] : x[91];
  assign t[169] = ~(t[176] & t[177]);
  assign t[16] = t[21] | t[22];
  assign t[170] = ~(t[272] & t[60]);
  assign t[171] = ~(t[277] & t[73]);
  assign t[172] = ~(t[284] & t[103]);
  assign t[173] = ~(t[287] & t[178]);
  assign t[174] = ~(t[274] & t[66]);
  assign t[175] = ~(t[91]);
  assign t[176] = ~(t[281] & t[96]);
  assign t[177] = ~(t[286] & t[179]);
  assign t[178] = ~(t[285] & t[102]);
  assign t[179] = ~(t[282] & t[95]);
  assign t[17] = ~(t[23] | t[24]);
  assign t[180] = t[1] ? t[181] : t[289];
  assign t[181] = x[6] ? t[183] : t[182];
  assign t[182] = x[7] ? t[185] : t[184];
  assign t[183] = t[186] ^ x[94];
  assign t[184] = t[187] ^ t[185];
  assign t[185] = ~(t[188] ^ t[189]);
  assign t[186] = x[95] ^ x[96];
  assign t[187] = t[262] ? x[95] : x[96];
  assign t[188] = x[7] ? t[191] : t[190];
  assign t[189] = ~(t[192] ^ t[193]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[190] = ~(t[194] & t[195]);
  assign t[191] = t[196] ^ t[197];
  assign t[192] = x[7] ? t[199] : t[198];
  assign t[193] = x[7] ? t[201] : t[200];
  assign t[194] = ~(t[36] & t[58]);
  assign t[195] = ~(t[202] & t[264]);
  assign t[196] = t[262] ? x[98] : x[97];
  assign t[197] = ~(t[203] & t[204]);
  assign t[198] = ~(t[205] & t[206]);
  assign t[199] = t[207] ^ t[208];
  assign t[19] = x[7] ? t[28] : t[27];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = ~(t[209] & t[210]);
  assign t[201] = t[211] ^ t[212];
  assign t[202] = ~(t[213] & t[35]);
  assign t[203] = ~(t[61] & t[89]);
  assign t[204] = ~(t[214] & t[267]);
  assign t[205] = ~(t[74] & t[100]);
  assign t[206] = ~(t[215] & t[269]);
  assign t[207] = t[262] ? x[100] : x[99];
  assign t[208] = ~(t[216] & t[217]);
  assign t[209] = ~(t[67] & t[93]);
  assign t[20] = x[7] ? t[30] : t[29];
  assign t[210] = ~(t[218] & t[268]);
  assign t[211] = t[219] ? x[102] : x[101];
  assign t[212] = ~(t[220] & t[221]);
  assign t[213] = ~(t[270] & t[266]);
  assign t[214] = ~(t[222] & t[60]);
  assign t[215] = ~(t[223] & t[73]);
  assign t[216] = ~(t[103] & t[119]);
  assign t[217] = ~(t[224] & t[278]);
  assign t[218] = ~(t[225] & t[66]);
  assign t[219] = ~(t[91]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = ~(t[96] & t[114]);
  assign t[221] = ~(t[226] & t[275]);
  assign t[222] = ~(t[279] & t[272]);
  assign t[223] = ~(t[283] & t[277]);
  assign t[224] = ~(t[227] & t[102]);
  assign t[225] = ~(t[280] & t[274]);
  assign t[226] = ~(t[228] & t[95]);
  assign t[227] = ~(t[287] & t[285]);
  assign t[228] = ~(t[286] & t[282]);
  assign t[229] = t[1] ? t[230] : t[290];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = x[6] ? t[232] : t[231];
  assign t[231] = x[7] ? t[234] : t[233];
  assign t[232] = t[235] ^ x[104];
  assign t[233] = t[236] ^ t[234];
  assign t[234] = ~(t[237] ^ t[238]);
  assign t[235] = x[105] ^ x[106];
  assign t[236] = t[262] ? x[105] : x[106];
  assign t[237] = x[7] ? t[240] : t[239];
  assign t[238] = ~(t[241] ^ t[242]);
  assign t[239] = ~(t[194] & t[243]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[240] = t[244] ^ t[245];
  assign t[241] = x[7] ? t[247] : t[246];
  assign t[242] = x[7] ? t[249] : t[248];
  assign t[243] = t[23] | t[264];
  assign t[244] = t[262] ? x[108] : x[107];
  assign t[245] = ~(t[203] & t[250]);
  assign t[246] = ~(t[205] & t[251]);
  assign t[247] = t[252] ^ t[253];
  assign t[248] = ~(t[209] & t[254]);
  assign t[249] = t[255] ^ t[256];
  assign t[24] = ~(t[264] | t[37]);
  assign t[250] = t[38] | t[267];
  assign t[251] = t[46] | t[269];
  assign t[252] = t[262] ? x[110] : x[109];
  assign t[253] = ~(t[216] & t[257]);
  assign t[254] = t[42] | t[268];
  assign t[255] = t[63] ? x[112] : x[111];
  assign t[256] = ~(t[220] & t[258]);
  assign t[257] = t[76] | t[278];
  assign t[258] = t[69] | t[275];
  assign t[259] = (t[291]);
  assign t[25] = ~(t[38] | t[39]);
  assign t[260] = (t[292]);
  assign t[261] = (t[293]);
  assign t[262] = (t[294]);
  assign t[263] = (t[295]);
  assign t[264] = (t[296]);
  assign t[265] = (t[297]);
  assign t[266] = (t[298]);
  assign t[267] = (t[299]);
  assign t[268] = (t[300]);
  assign t[269] = (t[301]);
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = (t[302]);
  assign t[271] = (t[303]);
  assign t[272] = (t[304]);
  assign t[273] = (t[305]);
  assign t[274] = (t[306]);
  assign t[275] = (t[307]);
  assign t[276] = (t[308]);
  assign t[277] = (t[309]);
  assign t[278] = (t[310]);
  assign t[279] = (t[311]);
  assign t[27] = ~(t[42] | t[43]);
  assign t[280] = (t[312]);
  assign t[281] = (t[313]);
  assign t[282] = (t[314]);
  assign t[283] = (t[315]);
  assign t[284] = (t[316]);
  assign t[285] = (t[317]);
  assign t[286] = (t[318]);
  assign t[287] = (t[319]);
  assign t[288] = (t[320]);
  assign t[289] = (t[321]);
  assign t[28] = ~(t[44] ^ t[45]);
  assign t[290] = (t[322]);
  assign t[291] = t[323] ^ x[5];
  assign t[292] = t[324] ^ x[11];
  assign t[293] = t[325] ^ x[14];
  assign t[294] = t[326] ^ x[17];
  assign t[295] = t[327] ^ x[20];
  assign t[296] = t[328] ^ x[28];
  assign t[297] = t[329] ^ x[29];
  assign t[298] = t[330] ^ x[30];
  assign t[299] = t[331] ^ x[36];
  assign t[29] = ~(t[46] | t[47]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = t[332] ^ x[44];
  assign t[301] = t[333] ^ x[50];
  assign t[302] = t[334] ^ x[51];
  assign t[303] = t[335] ^ x[52];
  assign t[304] = t[336] ^ x[53];
  assign t[305] = t[337] ^ x[54];
  assign t[306] = t[338] ^ x[55];
  assign t[307] = t[339] ^ x[61];
  assign t[308] = t[340] ^ x[64];
  assign t[309] = t[341] ^ x[65];
  assign t[30] = ~(t[48] ^ t[49]);
  assign t[310] = t[342] ^ x[71];
  assign t[311] = t[343] ^ x[74];
  assign t[312] = t[344] ^ x[75];
  assign t[313] = t[345] ^ x[76];
  assign t[314] = t[346] ^ x[77];
  assign t[315] = t[347] ^ x[78];
  assign t[316] = t[348] ^ x[79];
  assign t[317] = t[349] ^ x[80];
  assign t[318] = t[350] ^ x[81];
  assign t[319] = t[351] ^ x[82];
  assign t[31] = ~(t[50] & t[51]);
  assign t[320] = t[352] ^ x[83];
  assign t[321] = t[353] ^ x[93];
  assign t[322] = t[354] ^ x[103];
  assign t[323] = (~t[355] & t[356]);
  assign t[324] = (~t[357] & t[358]);
  assign t[325] = (~t[359] & t[360]);
  assign t[326] = (~t[361] & t[362]);
  assign t[327] = (~t[363] & t[364]);
  assign t[328] = (~t[365] & t[366]);
  assign t[329] = (~t[365] & t[367]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[330] = (~t[365] & t[368]);
  assign t[331] = (~t[369] & t[370]);
  assign t[332] = (~t[371] & t[372]);
  assign t[333] = (~t[373] & t[374]);
  assign t[334] = (~t[365] & t[375]);
  assign t[335] = (~t[369] & t[376]);
  assign t[336] = (~t[369] & t[377]);
  assign t[337] = (~t[371] & t[378]);
  assign t[338] = (~t[371] & t[379]);
  assign t[339] = (~t[380] & t[381]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = (~t[373] & t[382]);
  assign t[341] = (~t[373] & t[383]);
  assign t[342] = (~t[384] & t[385]);
  assign t[343] = (~t[369] & t[386]);
  assign t[344] = (~t[371] & t[387]);
  assign t[345] = (~t[380] & t[388]);
  assign t[346] = (~t[380] & t[389]);
  assign t[347] = (~t[373] & t[390]);
  assign t[348] = (~t[384] & t[391]);
  assign t[349] = (~t[384] & t[392]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[350] = (~t[380] & t[393]);
  assign t[351] = (~t[384] & t[394]);
  assign t[352] = (~t[355] & t[395]);
  assign t[353] = (~t[355] & t[396]);
  assign t[354] = (~t[355] & t[397]);
  assign t[355] = t[398] ^ x[4];
  assign t[356] = t[399] ^ x[5];
  assign t[357] = t[400] ^ x[10];
  assign t[358] = t[401] ^ x[11];
  assign t[359] = t[402] ^ x[13];
  assign t[35] = ~(t[265]);
  assign t[360] = t[403] ^ x[14];
  assign t[361] = t[404] ^ x[16];
  assign t[362] = t[405] ^ x[17];
  assign t[363] = t[406] ^ x[19];
  assign t[364] = t[407] ^ x[20];
  assign t[365] = t[408] ^ x[27];
  assign t[366] = t[409] ^ x[28];
  assign t[367] = t[410] ^ x[29];
  assign t[368] = t[411] ^ x[30];
  assign t[369] = t[412] ^ x[35];
  assign t[36] = ~(t[266]);
  assign t[370] = t[413] ^ x[36];
  assign t[371] = t[414] ^ x[43];
  assign t[372] = t[415] ^ x[44];
  assign t[373] = t[416] ^ x[49];
  assign t[374] = t[417] ^ x[50];
  assign t[375] = t[418] ^ x[51];
  assign t[376] = t[419] ^ x[52];
  assign t[377] = t[420] ^ x[53];
  assign t[378] = t[421] ^ x[54];
  assign t[379] = t[422] ^ x[55];
  assign t[37] = ~(t[58] | t[59]);
  assign t[380] = t[423] ^ x[60];
  assign t[381] = t[424] ^ x[61];
  assign t[382] = t[425] ^ x[64];
  assign t[383] = t[426] ^ x[65];
  assign t[384] = t[427] ^ x[70];
  assign t[385] = t[428] ^ x[71];
  assign t[386] = t[429] ^ x[74];
  assign t[387] = t[430] ^ x[75];
  assign t[388] = t[431] ^ x[76];
  assign t[389] = t[432] ^ x[77];
  assign t[38] = ~(t[60] | t[61]);
  assign t[390] = t[433] ^ x[78];
  assign t[391] = t[434] ^ x[79];
  assign t[392] = t[435] ^ x[80];
  assign t[393] = t[436] ^ x[81];
  assign t[394] = t[437] ^ x[82];
  assign t[395] = t[438] ^ x[83];
  assign t[396] = t[439] ^ x[93];
  assign t[397] = t[440] ^ x[103];
  assign t[398] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[399] = (x[0]);
  assign t[39] = ~(t[267] | t[62]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[401] = (x[9]);
  assign t[402] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[403] = (x[12]);
  assign t[404] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[405] = (x[15]);
  assign t[406] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[407] = (x[18]);
  assign t[408] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[409] = (x[24]);
  assign t[40] = t[63] ? x[38] : x[37];
  assign t[410] = (x[25]);
  assign t[411] = (x[26]);
  assign t[412] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[413] = (x[32]);
  assign t[414] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[415] = (x[40]);
  assign t[416] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[417] = (x[46]);
  assign t[418] = (x[23]);
  assign t[419] = (x[33]);
  assign t[41] = ~(t[64] & t[65]);
  assign t[420] = (x[34]);
  assign t[421] = (x[41]);
  assign t[422] = (x[42]);
  assign t[423] = (x[56] & ~x[57] & ~x[58] & ~x[59]) | (~x[56] & x[57] & ~x[58] & ~x[59]) | (~x[56] & ~x[57] & x[58] & ~x[59]) | (~x[56] & ~x[57] & ~x[58] & x[59]) | (x[56] & x[57] & x[58] & ~x[59]) | (x[56] & x[57] & ~x[58] & x[59]) | (x[56] & ~x[57] & x[58] & x[59]) | (~x[56] & x[57] & x[58] & x[59]);
  assign t[424] = (x[57]);
  assign t[425] = (x[47]);
  assign t[426] = (x[48]);
  assign t[427] = (x[66] & ~x[67] & ~x[68] & ~x[69]) | (~x[66] & x[67] & ~x[68] & ~x[69]) | (~x[66] & ~x[67] & x[68] & ~x[69]) | (~x[66] & ~x[67] & ~x[68] & x[69]) | (x[66] & x[67] & x[68] & ~x[69]) | (x[66] & x[67] & ~x[68] & x[69]) | (x[66] & ~x[67] & x[68] & x[69]) | (~x[66] & x[67] & x[68] & x[69]);
  assign t[428] = (x[67]);
  assign t[429] = (x[31]);
  assign t[42] = ~(t[66] | t[67]);
  assign t[430] = (x[39]);
  assign t[431] = (x[58]);
  assign t[432] = (x[59]);
  assign t[433] = (x[45]);
  assign t[434] = (x[68]);
  assign t[435] = (x[69]);
  assign t[436] = (x[56]);
  assign t[437] = (x[66]);
  assign t[438] = (x[1]);
  assign t[439] = (x[2]);
  assign t[43] = ~(t[268] | t[68]);
  assign t[440] = (x[3]);
  assign t[44] = ~(t[69] | t[70]);
  assign t[45] = ~(t[71] ^ t[72]);
  assign t[46] = ~(t[73] | t[74]);
  assign t[47] = ~(t[269] | t[75]);
  assign t[48] = ~(t[76] | t[77]);
  assign t[49] = ~(t[78] ^ t[79]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[80] | t[260]);
  assign t[51] = ~(t[81] & t[82]);
  assign t[52] = ~(t[261] | t[83]);
  assign t[53] = t[84] & t[260];
  assign t[54] = ~(t[84] | t[85]);
  assign t[55] = ~(t[84] | t[86]);
  assign t[56] = ~(t[84] | t[87]);
  assign t[57] = ~(t[84] | t[88]);
  assign t[58] = ~(t[270]);
  assign t[59] = ~(t[265] | t[266]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[271]);
  assign t[61] = ~(t[272]);
  assign t[62] = ~(t[89] | t[90]);
  assign t[63] = ~(t[91]);
  assign t[64] = ~(t[21] | t[92]);
  assign t[65] = ~(t[54]);
  assign t[66] = ~(t[273]);
  assign t[67] = ~(t[274]);
  assign t[68] = ~(t[93] | t[94]);
  assign t[69] = ~(t[95] | t[96]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[275] | t[97]);
  assign t[71] = t[262] ? x[63] : x[62];
  assign t[72] = ~(t[98] & t[99]);
  assign t[73] = ~(t[276]);
  assign t[74] = ~(t[277]);
  assign t[75] = ~(t[100] | t[101]);
  assign t[76] = ~(t[102] | t[103]);
  assign t[77] = ~(t[278] | t[104]);
  assign t[78] = t[262] ? x[73] : x[72];
  assign t[79] = ~(t[98] & t[105]);
  assign t[7] = ~(t[260] & t[261]);
  assign t[80] = ~(t[262]);
  assign t[81] = ~(t[263] & t[106]);
  assign t[82] = ~(x[7] & t[52]);
  assign t[83] = ~(t[263]);
  assign t[84] = ~(t[80]);
  assign t[85] = t[260] ? t[108] : t[107];
  assign t[86] = t[260] ? t[110] : t[109];
  assign t[87] = t[260] ? t[111] : t[81];
  assign t[88] = t[260] ? t[109] : t[110];
  assign t[89] = ~(t[279]);
  assign t[8] = ~(t[262] & t[263]);
  assign t[90] = ~(t[271] | t[272]);
  assign t[91] = ~(t[262]);
  assign t[92] = ~(t[112] & t[113]);
  assign t[93] = ~(t[280]);
  assign t[94] = ~(t[273] | t[274]);
  assign t[95] = ~(t[281]);
  assign t[96] = ~(t[282]);
  assign t[97] = ~(t[114] | t[115]);
  assign t[98] = ~(t[54] | t[116]);
  assign t[99] = ~(t[117] | t[118]);
  assign t[9] = ~(t[10] ^ t[12]);
  assign y = (t[0] & ~t[137] & ~t[180] & ~t[229]) | (~t[0] & t[137] & ~t[180] & ~t[229]) | (~t[0] & ~t[137] & t[180] & ~t[229]) | (~t[0] & ~t[137] & ~t[180] & t[229]) | (t[0] & t[137] & t[180] & ~t[229]) | (t[0] & t[137] & ~t[180] & t[229]) | (t[0] & ~t[137] & t[180] & t[229]) | (~t[0] & t[137] & t[180] & t[229]);
endmodule

module R2ind121(x, y);
 input [82:0] x;
 output y;

 wire [233:0] t;
  assign t[0] = t[1] ? t[2] : t[67];
  assign t[100] = t[129] ^ x[20];
  assign t[101] = t[130] ^ x[28];
  assign t[102] = t[131] ^ x[31];
  assign t[103] = t[132] ^ x[32];
  assign t[104] = t[133] ^ x[38];
  assign t[105] = t[134] ^ x[44];
  assign t[106] = t[135] ^ x[52];
  assign t[107] = t[136] ^ x[55];
  assign t[108] = t[137] ^ x[56];
  assign t[109] = t[138] ^ x[57];
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = t[139] ^ x[58];
  assign t[111] = t[140] ^ x[59];
  assign t[112] = t[141] ^ x[65];
  assign t[113] = t[142] ^ x[66];
  assign t[114] = t[143] ^ x[67];
  assign t[115] = t[144] ^ x[73];
  assign t[116] = t[145] ^ x[74];
  assign t[117] = t[146] ^ x[75];
  assign t[118] = t[147] ^ x[76];
  assign t[119] = t[148] ^ x[77];
  assign t[11] = x[21] ^ x[22];
  assign t[120] = t[149] ^ x[78];
  assign t[121] = t[150] ^ x[79];
  assign t[122] = t[151] ^ x[80];
  assign t[123] = t[152] ^ x[81];
  assign t[124] = t[153] ^ x[82];
  assign t[125] = (~t[154] & t[155]);
  assign t[126] = (~t[156] & t[157]);
  assign t[127] = (~t[158] & t[159]);
  assign t[128] = (~t[160] & t[161]);
  assign t[129] = (~t[162] & t[163]);
  assign t[12] = t[70] ? x[21] : x[22];
  assign t[130] = (~t[164] & t[165]);
  assign t[131] = (~t[164] & t[166]);
  assign t[132] = (~t[164] & t[167]);
  assign t[133] = (~t[168] & t[169]);
  assign t[134] = (~t[170] & t[171]);
  assign t[135] = (~t[172] & t[173]);
  assign t[136] = (~t[164] & t[174]);
  assign t[137] = (~t[168] & t[175]);
  assign t[138] = (~t[168] & t[176]);
  assign t[139] = (~t[170] & t[177]);
  assign t[13] = x[7] ? t[16] : t[15];
  assign t[140] = (~t[170] & t[178]);
  assign t[141] = (~t[179] & t[180]);
  assign t[142] = (~t[172] & t[181]);
  assign t[143] = (~t[172] & t[182]);
  assign t[144] = (~t[183] & t[184]);
  assign t[145] = (~t[168] & t[185]);
  assign t[146] = (~t[170] & t[186]);
  assign t[147] = (~t[179] & t[187]);
  assign t[148] = (~t[179] & t[188]);
  assign t[149] = (~t[172] & t[189]);
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = (~t[183] & t[190]);
  assign t[151] = (~t[183] & t[191]);
  assign t[152] = (~t[179] & t[192]);
  assign t[153] = (~t[183] & t[193]);
  assign t[154] = t[194] ^ x[4];
  assign t[155] = t[195] ^ x[5];
  assign t[156] = t[196] ^ x[10];
  assign t[157] = t[197] ^ x[11];
  assign t[158] = t[198] ^ x[13];
  assign t[159] = t[199] ^ x[14];
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[200] ^ x[16];
  assign t[161] = t[201] ^ x[17];
  assign t[162] = t[202] ^ x[19];
  assign t[163] = t[203] ^ x[20];
  assign t[164] = t[204] ^ x[27];
  assign t[165] = t[205] ^ x[28];
  assign t[166] = t[206] ^ x[31];
  assign t[167] = t[207] ^ x[32];
  assign t[168] = t[208] ^ x[37];
  assign t[169] = t[209] ^ x[38];
  assign t[16] = t[21] ^ t[22];
  assign t[170] = t[210] ^ x[43];
  assign t[171] = t[211] ^ x[44];
  assign t[172] = t[212] ^ x[51];
  assign t[173] = t[213] ^ x[52];
  assign t[174] = t[214] ^ x[55];
  assign t[175] = t[215] ^ x[56];
  assign t[176] = t[216] ^ x[57];
  assign t[177] = t[217] ^ x[58];
  assign t[178] = t[218] ^ x[59];
  assign t[179] = t[219] ^ x[64];
  assign t[17] = x[7] ? t[24] : t[23];
  assign t[180] = t[220] ^ x[65];
  assign t[181] = t[221] ^ x[66];
  assign t[182] = t[222] ^ x[67];
  assign t[183] = t[223] ^ x[72];
  assign t[184] = t[224] ^ x[73];
  assign t[185] = t[225] ^ x[74];
  assign t[186] = t[226] ^ x[75];
  assign t[187] = t[227] ^ x[76];
  assign t[188] = t[228] ^ x[77];
  assign t[189] = t[229] ^ x[78];
  assign t[18] = x[7] ? t[26] : t[25];
  assign t[190] = t[230] ^ x[79];
  assign t[191] = t[231] ^ x[80];
  assign t[192] = t[232] ^ x[81];
  assign t[193] = t[233] ^ x[82];
  assign t[194] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[195] = (x[3]);
  assign t[196] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[197] = (x[9]);
  assign t[198] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[199] = (x[12]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[201] = (x[15]);
  assign t[202] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[203] = (x[18]);
  assign t[204] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[205] = (x[24]);
  assign t[206] = (x[26]);
  assign t[207] = (x[23]);
  assign t[208] = (x[33] & ~x[34] & ~x[35] & ~x[36]) | (~x[33] & x[34] & ~x[35] & ~x[36]) | (~x[33] & ~x[34] & x[35] & ~x[36]) | (~x[33] & ~x[34] & ~x[35] & x[36]) | (x[33] & x[34] & x[35] & ~x[36]) | (x[33] & x[34] & ~x[35] & x[36]) | (x[33] & ~x[34] & x[35] & x[36]) | (~x[33] & x[34] & x[35] & x[36]);
  assign t[209] = (x[34]);
  assign t[20] = t[29] | t[72];
  assign t[210] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[211] = (x[40]);
  assign t[212] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[213] = (x[48]);
  assign t[214] = (x[25]);
  assign t[215] = (x[36]);
  assign t[216] = (x[33]);
  assign t[217] = (x[42]);
  assign t[218] = (x[39]);
  assign t[219] = (x[60] & ~x[61] & ~x[62] & ~x[63]) | (~x[60] & x[61] & ~x[62] & ~x[63]) | (~x[60] & ~x[61] & x[62] & ~x[63]) | (~x[60] & ~x[61] & ~x[62] & x[63]) | (x[60] & x[61] & x[62] & ~x[63]) | (x[60] & x[61] & ~x[62] & x[63]) | (x[60] & ~x[61] & x[62] & x[63]) | (~x[60] & x[61] & x[62] & x[63]);
  assign t[21] = t[70] ? x[30] : x[29];
  assign t[220] = (x[61]);
  assign t[221] = (x[50]);
  assign t[222] = (x[47]);
  assign t[223] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[224] = (x[69]);
  assign t[225] = (x[35]);
  assign t[226] = (x[41]);
  assign t[227] = (x[63]);
  assign t[228] = (x[60]);
  assign t[229] = (x[49]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[230] = (x[71]);
  assign t[231] = (x[68]);
  assign t[232] = (x[62]);
  assign t[233] = (x[70]);
  assign t[23] = ~(t[32] & t[33]);
  assign t[24] = t[34] ^ t[35];
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = ~(t[73]);
  assign t[28] = ~(t[74]);
  assign t[29] = ~(t[40] | t[27]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = ~(t[41] & t[42]);
  assign t[31] = t[43] | t[75];
  assign t[32] = ~(t[44] & t[45]);
  assign t[33] = t[46] | t[76];
  assign t[34] = t[70] ? x[46] : x[45];
  assign t[35] = ~(t[47] & t[48]);
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = t[51] | t[77];
  assign t[38] = t[52] ? x[54] : x[53];
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[78]);
  assign t[41] = ~(t[79]);
  assign t[42] = ~(t[80]);
  assign t[43] = ~(t[55] | t[41]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[82]);
  assign t[46] = ~(t[56] | t[44]);
  assign t[47] = ~(t[57] & t[58]);
  assign t[48] = t[59] | t[83];
  assign t[49] = ~(t[84]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[85]);
  assign t[51] = ~(t[60] | t[49]);
  assign t[52] = ~(t[61]);
  assign t[53] = ~(t[62] & t[63]);
  assign t[54] = t[64] | t[86];
  assign t[55] = ~(t[87]);
  assign t[56] = ~(t[88]);
  assign t[57] = ~(t[89]);
  assign t[58] = ~(t[90]);
  assign t[59] = ~(t[65] | t[57]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[91]);
  assign t[61] = ~(t[70]);
  assign t[62] = ~(t[92]);
  assign t[63] = ~(t[93]);
  assign t[64] = ~(t[66] | t[62]);
  assign t[65] = ~(t[94]);
  assign t[66] = ~(t[95]);
  assign t[67] = (t[96]);
  assign t[68] = (t[97]);
  assign t[69] = (t[98]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = (t[99]);
  assign t[71] = (t[100]);
  assign t[72] = (t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = ~(t[68] & t[69]);
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[70] & t[71]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = t[125] ^ x[5];
  assign t[97] = t[126] ^ x[11];
  assign t[98] = t[127] ^ x[14];
  assign t[99] = t[128] ^ x[17];
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [82:0] x;
 output y;

 wire [239:0] t;
  assign t[0] = t[1] ? t[2] : t[73];
  assign t[100] = (t[129]);
  assign t[101] = (t[130]);
  assign t[102] = t[131] ^ x[5];
  assign t[103] = t[132] ^ x[11];
  assign t[104] = t[133] ^ x[14];
  assign t[105] = t[134] ^ x[17];
  assign t[106] = t[135] ^ x[20];
  assign t[107] = t[136] ^ x[28];
  assign t[108] = t[137] ^ x[31];
  assign t[109] = t[138] ^ x[32];
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = t[139] ^ x[38];
  assign t[111] = t[140] ^ x[44];
  assign t[112] = t[141] ^ x[52];
  assign t[113] = t[142] ^ x[55];
  assign t[114] = t[143] ^ x[56];
  assign t[115] = t[144] ^ x[57];
  assign t[116] = t[145] ^ x[58];
  assign t[117] = t[146] ^ x[59];
  assign t[118] = t[147] ^ x[65];
  assign t[119] = t[148] ^ x[66];
  assign t[11] = x[21] ^ x[22];
  assign t[120] = t[149] ^ x[67];
  assign t[121] = t[150] ^ x[73];
  assign t[122] = t[151] ^ x[74];
  assign t[123] = t[152] ^ x[75];
  assign t[124] = t[153] ^ x[76];
  assign t[125] = t[154] ^ x[77];
  assign t[126] = t[155] ^ x[78];
  assign t[127] = t[156] ^ x[79];
  assign t[128] = t[157] ^ x[80];
  assign t[129] = t[158] ^ x[81];
  assign t[12] = t[76] ? x[21] : x[22];
  assign t[130] = t[159] ^ x[82];
  assign t[131] = (~t[160] & t[161]);
  assign t[132] = (~t[162] & t[163]);
  assign t[133] = (~t[164] & t[165]);
  assign t[134] = (~t[166] & t[167]);
  assign t[135] = (~t[168] & t[169]);
  assign t[136] = (~t[170] & t[171]);
  assign t[137] = (~t[170] & t[172]);
  assign t[138] = (~t[170] & t[173]);
  assign t[139] = (~t[174] & t[175]);
  assign t[13] = x[7] ? t[16] : t[15];
  assign t[140] = (~t[176] & t[177]);
  assign t[141] = (~t[178] & t[179]);
  assign t[142] = (~t[170] & t[180]);
  assign t[143] = (~t[174] & t[181]);
  assign t[144] = (~t[174] & t[182]);
  assign t[145] = (~t[176] & t[183]);
  assign t[146] = (~t[176] & t[184]);
  assign t[147] = (~t[185] & t[186]);
  assign t[148] = (~t[178] & t[187]);
  assign t[149] = (~t[178] & t[188]);
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = (~t[189] & t[190]);
  assign t[151] = (~t[174] & t[191]);
  assign t[152] = (~t[176] & t[192]);
  assign t[153] = (~t[185] & t[193]);
  assign t[154] = (~t[185] & t[194]);
  assign t[155] = (~t[178] & t[195]);
  assign t[156] = (~t[189] & t[196]);
  assign t[157] = (~t[189] & t[197]);
  assign t[158] = (~t[185] & t[198]);
  assign t[159] = (~t[189] & t[199]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[200] ^ x[4];
  assign t[161] = t[201] ^ x[5];
  assign t[162] = t[202] ^ x[10];
  assign t[163] = t[203] ^ x[11];
  assign t[164] = t[204] ^ x[13];
  assign t[165] = t[205] ^ x[14];
  assign t[166] = t[206] ^ x[16];
  assign t[167] = t[207] ^ x[17];
  assign t[168] = t[208] ^ x[19];
  assign t[169] = t[209] ^ x[20];
  assign t[16] = t[21] ^ t[22];
  assign t[170] = t[210] ^ x[27];
  assign t[171] = t[211] ^ x[28];
  assign t[172] = t[212] ^ x[31];
  assign t[173] = t[213] ^ x[32];
  assign t[174] = t[214] ^ x[37];
  assign t[175] = t[215] ^ x[38];
  assign t[176] = t[216] ^ x[43];
  assign t[177] = t[217] ^ x[44];
  assign t[178] = t[218] ^ x[51];
  assign t[179] = t[219] ^ x[52];
  assign t[17] = x[7] ? t[24] : t[23];
  assign t[180] = t[220] ^ x[55];
  assign t[181] = t[221] ^ x[56];
  assign t[182] = t[222] ^ x[57];
  assign t[183] = t[223] ^ x[58];
  assign t[184] = t[224] ^ x[59];
  assign t[185] = t[225] ^ x[64];
  assign t[186] = t[226] ^ x[65];
  assign t[187] = t[227] ^ x[66];
  assign t[188] = t[228] ^ x[67];
  assign t[189] = t[229] ^ x[72];
  assign t[18] = x[7] ? t[26] : t[25];
  assign t[190] = t[230] ^ x[73];
  assign t[191] = t[231] ^ x[74];
  assign t[192] = t[232] ^ x[75];
  assign t[193] = t[233] ^ x[76];
  assign t[194] = t[234] ^ x[77];
  assign t[195] = t[235] ^ x[78];
  assign t[196] = t[236] ^ x[79];
  assign t[197] = t[237] ^ x[80];
  assign t[198] = t[238] ^ x[81];
  assign t[199] = t[239] ^ x[82];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[201] = (x[2]);
  assign t[202] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[203] = (x[9]);
  assign t[204] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[205] = (x[12]);
  assign t[206] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[207] = (x[15]);
  assign t[208] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[209] = (x[18]);
  assign t[20] = ~(t[29] & t[78]);
  assign t[210] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[211] = (x[24]);
  assign t[212] = (x[26]);
  assign t[213] = (x[23]);
  assign t[214] = (x[33] & ~x[34] & ~x[35] & ~x[36]) | (~x[33] & x[34] & ~x[35] & ~x[36]) | (~x[33] & ~x[34] & x[35] & ~x[36]) | (~x[33] & ~x[34] & ~x[35] & x[36]) | (x[33] & x[34] & x[35] & ~x[36]) | (x[33] & x[34] & ~x[35] & x[36]) | (x[33] & ~x[34] & x[35] & x[36]) | (~x[33] & x[34] & x[35] & x[36]);
  assign t[215] = (x[34]);
  assign t[216] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[217] = (x[40]);
  assign t[218] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[219] = (x[48]);
  assign t[21] = t[76] ? x[30] : x[29];
  assign t[220] = (x[25]);
  assign t[221] = (x[36]);
  assign t[222] = (x[33]);
  assign t[223] = (x[42]);
  assign t[224] = (x[39]);
  assign t[225] = (x[60] & ~x[61] & ~x[62] & ~x[63]) | (~x[60] & x[61] & ~x[62] & ~x[63]) | (~x[60] & ~x[61] & x[62] & ~x[63]) | (~x[60] & ~x[61] & ~x[62] & x[63]) | (x[60] & x[61] & x[62] & ~x[63]) | (x[60] & x[61] & ~x[62] & x[63]) | (x[60] & ~x[61] & x[62] & x[63]) | (~x[60] & x[61] & x[62] & x[63]);
  assign t[226] = (x[61]);
  assign t[227] = (x[50]);
  assign t[228] = (x[47]);
  assign t[229] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[230] = (x[69]);
  assign t[231] = (x[35]);
  assign t[232] = (x[41]);
  assign t[233] = (x[63]);
  assign t[234] = (x[60]);
  assign t[235] = (x[49]);
  assign t[236] = (x[71]);
  assign t[237] = (x[68]);
  assign t[238] = (x[62]);
  assign t[239] = (x[70]);
  assign t[23] = ~(t[32] & t[33]);
  assign t[24] = t[34] ^ t[35];
  assign t[25] = ~(t[36] & t[37]);
  assign t[26] = t[38] ^ t[39];
  assign t[27] = ~(t[79]);
  assign t[28] = ~(t[80]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = ~(t[42] & t[43]);
  assign t[31] = ~(t[44] & t[81]);
  assign t[32] = ~(t[45] & t[46]);
  assign t[33] = ~(t[47] & t[82]);
  assign t[34] = t[76] ? x[46] : x[45];
  assign t[35] = ~(t[48] & t[49]);
  assign t[36] = ~(t[50] & t[51]);
  assign t[37] = ~(t[52] & t[83]);
  assign t[38] = t[53] ? x[54] : x[53];
  assign t[39] = ~(t[54] & t[55]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[80] & t[79]);
  assign t[41] = ~(t[84]);
  assign t[42] = ~(t[85]);
  assign t[43] = ~(t[86]);
  assign t[44] = ~(t[56] & t[57]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[88]);
  assign t[47] = ~(t[58] & t[59]);
  assign t[48] = ~(t[60] & t[61]);
  assign t[49] = ~(t[62] & t[89]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[90]);
  assign t[51] = ~(t[91]);
  assign t[52] = ~(t[63] & t[64]);
  assign t[53] = ~(t[65]);
  assign t[54] = ~(t[66] & t[67]);
  assign t[55] = ~(t[68] & t[92]);
  assign t[56] = ~(t[86] & t[85]);
  assign t[57] = ~(t[93]);
  assign t[58] = ~(t[88] & t[87]);
  assign t[59] = ~(t[94]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[95]);
  assign t[61] = ~(t[96]);
  assign t[62] = ~(t[69] & t[70]);
  assign t[63] = ~(t[91] & t[90]);
  assign t[64] = ~(t[97]);
  assign t[65] = ~(t[76]);
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[99]);
  assign t[68] = ~(t[71] & t[72]);
  assign t[69] = ~(t[96] & t[95]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[100]);
  assign t[71] = ~(t[99] & t[98]);
  assign t[72] = ~(t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = ~(t[74] & t[75]);
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[76] & t[77]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = (t[128]);
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [76:0] x;
 output y;

 wire [197:0] t;
  assign t[0] = t[1] ? t[2] : t[61];
  assign t[100] = t[123] ^ x[65];
  assign t[101] = t[124] ^ x[66];
  assign t[102] = t[125] ^ x[67];
  assign t[103] = t[126] ^ x[73];
  assign t[104] = t[127] ^ x[74];
  assign t[105] = t[128] ^ x[75];
  assign t[106] = t[129] ^ x[76];
  assign t[107] = (~t[130] & t[131]);
  assign t[108] = (~t[132] & t[133]);
  assign t[109] = (~t[134] & t[135]);
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = (~t[136] & t[137]);
  assign t[111] = (~t[138] & t[139]);
  assign t[112] = (~t[140] & t[141]);
  assign t[113] = (~t[140] & t[142]);
  assign t[114] = (~t[140] & t[143]);
  assign t[115] = (~t[144] & t[145]);
  assign t[116] = (~t[144] & t[146]);
  assign t[117] = (~t[147] & t[148]);
  assign t[118] = (~t[147] & t[149]);
  assign t[119] = (~t[150] & t[151]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (~t[150] & t[152]);
  assign t[121] = (~t[144] & t[153]);
  assign t[122] = (~t[147] & t[154]);
  assign t[123] = (~t[155] & t[156]);
  assign t[124] = (~t[155] & t[157]);
  assign t[125] = (~t[150] & t[158]);
  assign t[126] = (~t[159] & t[160]);
  assign t[127] = (~t[159] & t[161]);
  assign t[128] = (~t[155] & t[162]);
  assign t[129] = (~t[159] & t[163]);
  assign t[12] = t[64] ? x[22] : x[21];
  assign t[130] = t[164] ^ x[4];
  assign t[131] = t[165] ^ x[5];
  assign t[132] = t[166] ^ x[10];
  assign t[133] = t[167] ^ x[11];
  assign t[134] = t[168] ^ x[13];
  assign t[135] = t[169] ^ x[14];
  assign t[136] = t[170] ^ x[16];
  assign t[137] = t[171] ^ x[17];
  assign t[138] = t[172] ^ x[19];
  assign t[139] = t[173] ^ x[20];
  assign t[13] = x[7] ? t[16] : t[15];
  assign t[140] = t[174] ^ x[27];
  assign t[141] = t[175] ^ x[28];
  assign t[142] = t[176] ^ x[29];
  assign t[143] = t[177] ^ x[32];
  assign t[144] = t[178] ^ x[37];
  assign t[145] = t[179] ^ x[38];
  assign t[146] = t[180] ^ x[39];
  assign t[147] = t[181] ^ x[44];
  assign t[148] = t[182] ^ x[45];
  assign t[149] = t[183] ^ x[46];
  assign t[14] = ~(t[17] ^ t[18]);
  assign t[150] = t[184] ^ x[53];
  assign t[151] = t[185] ^ x[54];
  assign t[152] = t[186] ^ x[55];
  assign t[153] = t[187] ^ x[58];
  assign t[154] = t[188] ^ x[59];
  assign t[155] = t[189] ^ x[64];
  assign t[156] = t[190] ^ x[65];
  assign t[157] = t[191] ^ x[66];
  assign t[158] = t[192] ^ x[67];
  assign t[159] = t[193] ^ x[72];
  assign t[15] = ~(t[19] & t[20]);
  assign t[160] = t[194] ^ x[73];
  assign t[161] = t[195] ^ x[74];
  assign t[162] = t[196] ^ x[75];
  assign t[163] = t[197] ^ x[76];
  assign t[164] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[165] = (x[1]);
  assign t[166] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[167] = (x[9]);
  assign t[168] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[169] = (x[12]);
  assign t[16] = t[21] ^ t[22];
  assign t[170] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[171] = (x[15]);
  assign t[172] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[173] = (x[18]);
  assign t[174] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[175] = (x[25]);
  assign t[176] = (x[23]);
  assign t[177] = (x[26]);
  assign t[178] = (x[33] & ~x[34] & ~x[35] & ~x[36]) | (~x[33] & x[34] & ~x[35] & ~x[36]) | (~x[33] & ~x[34] & x[35] & ~x[36]) | (~x[33] & ~x[34] & ~x[35] & x[36]) | (x[33] & x[34] & x[35] & ~x[36]) | (x[33] & x[34] & ~x[35] & x[36]) | (x[33] & ~x[34] & x[35] & x[36]) | (~x[33] & x[34] & x[35] & x[36]);
  assign t[179] = (x[35]);
  assign t[17] = x[7] ? t[24] : t[23];
  assign t[180] = (x[33]);
  assign t[181] = (x[40] & ~x[41] & ~x[42] & ~x[43]) | (~x[40] & x[41] & ~x[42] & ~x[43]) | (~x[40] & ~x[41] & x[42] & ~x[43]) | (~x[40] & ~x[41] & ~x[42] & x[43]) | (x[40] & x[41] & x[42] & ~x[43]) | (x[40] & x[41] & ~x[42] & x[43]) | (x[40] & ~x[41] & x[42] & x[43]) | (~x[40] & x[41] & x[42] & x[43]);
  assign t[182] = (x[42]);
  assign t[183] = (x[40]);
  assign t[184] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[185] = (x[51]);
  assign t[186] = (x[49]);
  assign t[187] = (x[36]);
  assign t[188] = (x[43]);
  assign t[189] = (x[60] & ~x[61] & ~x[62] & ~x[63]) | (~x[60] & x[61] & ~x[62] & ~x[63]) | (~x[60] & ~x[61] & x[62] & ~x[63]) | (~x[60] & ~x[61] & ~x[62] & x[63]) | (x[60] & x[61] & x[62] & ~x[63]) | (x[60] & x[61] & ~x[62] & x[63]) | (x[60] & ~x[61] & x[62] & x[63]) | (~x[60] & x[61] & x[62] & x[63]);
  assign t[18] = x[7] ? t[26] : t[25];
  assign t[190] = (x[62]);
  assign t[191] = (x[60]);
  assign t[192] = (x[52]);
  assign t[193] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[194] = (x[70]);
  assign t[195] = (x[68]);
  assign t[196] = (x[63]);
  assign t[197] = (x[71]);
  assign t[19] = ~(t[66] & t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[67] & t[28]);
  assign t[21] = t[64] ? x[31] : x[30];
  assign t[22] = ~(t[29] & t[30]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[35] & t[36]);
  assign t[26] = t[37] ^ t[38];
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[68] & t[39]);
  assign t[29] = ~(t[69] & t[40]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = ~(t[70] & t[41]);
  assign t[31] = ~(t[71] & t[42]);
  assign t[32] = ~(t[72] & t[43]);
  assign t[33] = t[64] ? x[48] : x[47];
  assign t[34] = ~(t[44] & t[45]);
  assign t[35] = ~(t[73] & t[46]);
  assign t[36] = ~(t[74] & t[47]);
  assign t[37] = t[48] ? x[57] : x[56];
  assign t[38] = ~(t[49] & t[50]);
  assign t[39] = ~(t[66]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[75]);
  assign t[41] = ~(t[75] & t[51]);
  assign t[42] = ~(t[76]);
  assign t[43] = ~(t[76] & t[52]);
  assign t[44] = ~(t[77] & t[53]);
  assign t[45] = ~(t[78] & t[54]);
  assign t[46] = ~(t[79]);
  assign t[47] = ~(t[79] & t[55]);
  assign t[48] = ~(t[56]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[81] & t[58]);
  assign t[51] = ~(t[69]);
  assign t[52] = ~(t[71]);
  assign t[53] = ~(t[82]);
  assign t[54] = ~(t[82] & t[59]);
  assign t[55] = ~(t[73]);
  assign t[56] = ~(t[64]);
  assign t[57] = ~(t[83]);
  assign t[58] = ~(t[83] & t[60]);
  assign t[59] = ~(t[77]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[80]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = (t[86]);
  assign t[64] = (t[87]);
  assign t[65] = (t[88]);
  assign t[66] = (t[89]);
  assign t[67] = (t[90]);
  assign t[68] = (t[91]);
  assign t[69] = (t[92]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = (t[93]);
  assign t[71] = (t[94]);
  assign t[72] = (t[95]);
  assign t[73] = (t[96]);
  assign t[74] = (t[97]);
  assign t[75] = (t[98]);
  assign t[76] = (t[99]);
  assign t[77] = (t[100]);
  assign t[78] = (t[101]);
  assign t[79] = (t[102]);
  assign t[7] = ~(t[62] & t[63]);
  assign t[80] = (t[103]);
  assign t[81] = (t[104]);
  assign t[82] = (t[105]);
  assign t[83] = (t[106]);
  assign t[84] = t[107] ^ x[5];
  assign t[85] = t[108] ^ x[11];
  assign t[86] = t[109] ^ x[14];
  assign t[87] = t[110] ^ x[17];
  assign t[88] = t[111] ^ x[20];
  assign t[89] = t[112] ^ x[28];
  assign t[8] = ~(t[64] & t[65]);
  assign t[90] = t[113] ^ x[29];
  assign t[91] = t[114] ^ x[32];
  assign t[92] = t[115] ^ x[38];
  assign t[93] = t[116] ^ x[39];
  assign t[94] = t[117] ^ x[45];
  assign t[95] = t[118] ^ x[46];
  assign t[96] = t[119] ^ x[54];
  assign t[97] = t[120] ^ x[55];
  assign t[98] = t[121] ^ x[58];
  assign t[99] = t[122] ^ x[59];
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [82:0] x;
 output y;

 wire [303:0] t;
  assign t[0] = t[1] ? t[2] : t[137];
  assign t[100] = ~(t[161]);
  assign t[101] = ~(t[154] | t[155]);
  assign t[102] = ~(t[162]);
  assign t[103] = ~(t[163]);
  assign t[104] = ~(t[119] | t[120]);
  assign t[105] = ~(t[121] | t[57]);
  assign t[106] = ~(x[7] | t[122]);
  assign t[107] = ~(t[123] & t[141]);
  assign t[108] = ~(t[124] & t[83]);
  assign t[109] = ~(t[123] & t[83]);
  assign t[10] = ~(t[13] ^ t[14]);
  assign t[110] = ~(t[124] & t[141]);
  assign t[111] = ~(x[7] & t[125]);
  assign t[112] = ~(t[117]);
  assign t[113] = t[80] | t[126];
  assign t[114] = ~(t[164]);
  assign t[115] = ~(t[159] | t[160]);
  assign t[116] = ~(t[127] & t[128]);
  assign t[117] = ~(t[80] | t[129]);
  assign t[118] = t[55] | t[130];
  assign t[119] = ~(t[165]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = ~(t[162] | t[163]);
  assign t[121] = ~(t[84] | t[131]);
  assign t[122] = ~(t[139]);
  assign t[123] = x[7] & t[139];
  assign t[124] = ~(x[7] | t[139]);
  assign t[125] = ~(t[139] | t[141]);
  assign t[126] = t[138] ? t[111] : t[132];
  assign t[127] = ~(t[133] | t[56]);
  assign t[128] = ~(t[134] & t[135]);
  assign t[129] = t[138] ? t[132] : t[111];
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[130] = ~(t[31]);
  assign t[131] = t[138] ? t[82] : t[132];
  assign t[132] = ~(t[106] & t[83]);
  assign t[133] = ~(t[84] | t[136]);
  assign t[134] = t[141] & t[50];
  assign t[135] = t[124] | t[123];
  assign t[136] = t[138] ? t[107] : t[108];
  assign t[137] = (t[166]);
  assign t[138] = (t[167]);
  assign t[139] = (t[168]);
  assign t[13] = x[7] ? t[18] : t[17];
  assign t[140] = (t[169]);
  assign t[141] = (t[170]);
  assign t[142] = (t[171]);
  assign t[143] = (t[172]);
  assign t[144] = (t[173]);
  assign t[145] = (t[174]);
  assign t[146] = (t[175]);
  assign t[147] = (t[176]);
  assign t[148] = (t[177]);
  assign t[149] = (t[178]);
  assign t[14] = ~(t[19] ^ t[20]);
  assign t[150] = (t[179]);
  assign t[151] = (t[180]);
  assign t[152] = (t[181]);
  assign t[153] = (t[182]);
  assign t[154] = (t[183]);
  assign t[155] = (t[184]);
  assign t[156] = (t[185]);
  assign t[157] = (t[186]);
  assign t[158] = (t[187]);
  assign t[159] = (t[188]);
  assign t[15] = t[140] ? x[22] : x[21];
  assign t[160] = (t[189]);
  assign t[161] = (t[190]);
  assign t[162] = (t[191]);
  assign t[163] = (t[192]);
  assign t[164] = (t[193]);
  assign t[165] = (t[194]);
  assign t[166] = t[195] ^ x[5];
  assign t[167] = t[196] ^ x[11];
  assign t[168] = t[197] ^ x[14];
  assign t[169] = t[198] ^ x[17];
  assign t[16] = t[21] | t[22];
  assign t[170] = t[199] ^ x[20];
  assign t[171] = t[200] ^ x[28];
  assign t[172] = t[201] ^ x[29];
  assign t[173] = t[202] ^ x[30];
  assign t[174] = t[203] ^ x[36];
  assign t[175] = t[204] ^ x[44];
  assign t[176] = t[205] ^ x[50];
  assign t[177] = t[206] ^ x[51];
  assign t[178] = t[207] ^ x[52];
  assign t[179] = t[208] ^ x[53];
  assign t[17] = ~(t[23] | t[24]);
  assign t[180] = t[209] ^ x[54];
  assign t[181] = t[210] ^ x[55];
  assign t[182] = t[211] ^ x[61];
  assign t[183] = t[212] ^ x[64];
  assign t[184] = t[213] ^ x[65];
  assign t[185] = t[214] ^ x[71];
  assign t[186] = t[215] ^ x[74];
  assign t[187] = t[216] ^ x[75];
  assign t[188] = t[217] ^ x[76];
  assign t[189] = t[218] ^ x[77];
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[190] = t[219] ^ x[78];
  assign t[191] = t[220] ^ x[79];
  assign t[192] = t[221] ^ x[80];
  assign t[193] = t[222] ^ x[81];
  assign t[194] = t[223] ^ x[82];
  assign t[195] = (~t[224] & t[225]);
  assign t[196] = (~t[226] & t[227]);
  assign t[197] = (~t[228] & t[229]);
  assign t[198] = (~t[230] & t[231]);
  assign t[199] = (~t[232] & t[233]);
  assign t[19] = x[7] ? t[28] : t[27];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (~t[234] & t[235]);
  assign t[201] = (~t[234] & t[236]);
  assign t[202] = (~t[234] & t[237]);
  assign t[203] = (~t[238] & t[239]);
  assign t[204] = (~t[240] & t[241]);
  assign t[205] = (~t[242] & t[243]);
  assign t[206] = (~t[234] & t[244]);
  assign t[207] = (~t[238] & t[245]);
  assign t[208] = (~t[238] & t[246]);
  assign t[209] = (~t[240] & t[247]);
  assign t[20] = x[7] ? t[30] : t[29];
  assign t[210] = (~t[240] & t[248]);
  assign t[211] = (~t[249] & t[250]);
  assign t[212] = (~t[242] & t[251]);
  assign t[213] = (~t[242] & t[252]);
  assign t[214] = (~t[253] & t[254]);
  assign t[215] = (~t[238] & t[255]);
  assign t[216] = (~t[240] & t[256]);
  assign t[217] = (~t[249] & t[257]);
  assign t[218] = (~t[249] & t[258]);
  assign t[219] = (~t[242] & t[259]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (~t[253] & t[260]);
  assign t[221] = (~t[253] & t[261]);
  assign t[222] = (~t[249] & t[262]);
  assign t[223] = (~t[253] & t[263]);
  assign t[224] = t[264] ^ x[4];
  assign t[225] = t[265] ^ x[5];
  assign t[226] = t[266] ^ x[10];
  assign t[227] = t[267] ^ x[11];
  assign t[228] = t[268] ^ x[13];
  assign t[229] = t[269] ^ x[14];
  assign t[22] = ~(t[33] & t[34]);
  assign t[230] = t[270] ^ x[16];
  assign t[231] = t[271] ^ x[17];
  assign t[232] = t[272] ^ x[19];
  assign t[233] = t[273] ^ x[20];
  assign t[234] = t[274] ^ x[27];
  assign t[235] = t[275] ^ x[28];
  assign t[236] = t[276] ^ x[29];
  assign t[237] = t[277] ^ x[30];
  assign t[238] = t[278] ^ x[35];
  assign t[239] = t[279] ^ x[36];
  assign t[23] = ~(t[35] | t[36]);
  assign t[240] = t[280] ^ x[43];
  assign t[241] = t[281] ^ x[44];
  assign t[242] = t[282] ^ x[49];
  assign t[243] = t[283] ^ x[50];
  assign t[244] = t[284] ^ x[51];
  assign t[245] = t[285] ^ x[52];
  assign t[246] = t[286] ^ x[53];
  assign t[247] = t[287] ^ x[54];
  assign t[248] = t[288] ^ x[55];
  assign t[249] = t[289] ^ x[60];
  assign t[24] = ~(t[142] | t[37]);
  assign t[250] = t[290] ^ x[61];
  assign t[251] = t[291] ^ x[64];
  assign t[252] = t[292] ^ x[65];
  assign t[253] = t[293] ^ x[70];
  assign t[254] = t[294] ^ x[71];
  assign t[255] = t[295] ^ x[74];
  assign t[256] = t[296] ^ x[75];
  assign t[257] = t[297] ^ x[76];
  assign t[258] = t[298] ^ x[77];
  assign t[259] = t[299] ^ x[78];
  assign t[25] = ~(t[38] | t[39]);
  assign t[260] = t[300] ^ x[79];
  assign t[261] = t[301] ^ x[80];
  assign t[262] = t[302] ^ x[81];
  assign t[263] = t[303] ^ x[82];
  assign t[264] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[265] = (x[0]);
  assign t[266] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[267] = (x[9]);
  assign t[268] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[269] = (x[12]);
  assign t[26] = ~(t[40] ^ t[41]);
  assign t[270] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[271] = (x[15]);
  assign t[272] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[273] = (x[18]);
  assign t[274] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[275] = (x[24]);
  assign t[276] = (x[25]);
  assign t[277] = (x[26]);
  assign t[278] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[279] = (x[32]);
  assign t[27] = ~(t[42] | t[43]);
  assign t[280] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[281] = (x[40]);
  assign t[282] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[283] = (x[46]);
  assign t[284] = (x[23]);
  assign t[285] = (x[33]);
  assign t[286] = (x[34]);
  assign t[287] = (x[41]);
  assign t[288] = (x[42]);
  assign t[289] = (x[56] & ~x[57] & ~x[58] & ~x[59]) | (~x[56] & x[57] & ~x[58] & ~x[59]) | (~x[56] & ~x[57] & x[58] & ~x[59]) | (~x[56] & ~x[57] & ~x[58] & x[59]) | (x[56] & x[57] & x[58] & ~x[59]) | (x[56] & x[57] & ~x[58] & x[59]) | (x[56] & ~x[57] & x[58] & x[59]) | (~x[56] & x[57] & x[58] & x[59]);
  assign t[28] = ~(t[44] ^ t[45]);
  assign t[290] = (x[57]);
  assign t[291] = (x[47]);
  assign t[292] = (x[48]);
  assign t[293] = (x[66] & ~x[67] & ~x[68] & ~x[69]) | (~x[66] & x[67] & ~x[68] & ~x[69]) | (~x[66] & ~x[67] & x[68] & ~x[69]) | (~x[66] & ~x[67] & ~x[68] & x[69]) | (x[66] & x[67] & x[68] & ~x[69]) | (x[66] & x[67] & ~x[68] & x[69]) | (x[66] & ~x[67] & x[68] & x[69]) | (~x[66] & x[67] & x[68] & x[69]);
  assign t[294] = (x[67]);
  assign t[295] = (x[31]);
  assign t[296] = (x[39]);
  assign t[297] = (x[58]);
  assign t[298] = (x[59]);
  assign t[299] = (x[45]);
  assign t[29] = ~(t[46] | t[47]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = (x[68]);
  assign t[301] = (x[69]);
  assign t[302] = (x[56]);
  assign t[303] = (x[66]);
  assign t[30] = ~(t[48] ^ t[49]);
  assign t[31] = ~(t[50] & t[51]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[34] = ~(t[56] | t[57]);
  assign t[35] = ~(t[143]);
  assign t[36] = ~(t[144]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = ~(t[60] | t[61]);
  assign t[39] = ~(t[145] | t[62]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[63] ? x[38] : x[37];
  assign t[41] = ~(t[64] & t[65]);
  assign t[42] = ~(t[66] | t[67]);
  assign t[43] = ~(t[146] | t[68]);
  assign t[44] = ~(t[69] | t[70]);
  assign t[45] = ~(t[71] ^ t[72]);
  assign t[46] = ~(t[73] | t[74]);
  assign t[47] = ~(t[147] | t[75]);
  assign t[48] = ~(t[76] | t[77]);
  assign t[49] = ~(t[78] ^ t[79]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[80] | t[138]);
  assign t[51] = ~(t[81] & t[82]);
  assign t[52] = ~(t[139] | t[83]);
  assign t[53] = t[84] & t[138];
  assign t[54] = ~(t[84] | t[85]);
  assign t[55] = ~(t[84] | t[86]);
  assign t[56] = ~(t[84] | t[87]);
  assign t[57] = ~(t[84] | t[88]);
  assign t[58] = ~(t[148]);
  assign t[59] = ~(t[143] | t[144]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[149]);
  assign t[61] = ~(t[150]);
  assign t[62] = ~(t[89] | t[90]);
  assign t[63] = ~(t[91]);
  assign t[64] = ~(t[21] | t[92]);
  assign t[65] = ~(t[54]);
  assign t[66] = ~(t[151]);
  assign t[67] = ~(t[152]);
  assign t[68] = ~(t[93] | t[94]);
  assign t[69] = ~(t[95] | t[96]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[153] | t[97]);
  assign t[71] = t[140] ? x[63] : x[62];
  assign t[72] = ~(t[98] & t[99]);
  assign t[73] = ~(t[154]);
  assign t[74] = ~(t[155]);
  assign t[75] = ~(t[100] | t[101]);
  assign t[76] = ~(t[102] | t[103]);
  assign t[77] = ~(t[156] | t[104]);
  assign t[78] = t[140] ? x[73] : x[72];
  assign t[79] = ~(t[98] & t[105]);
  assign t[7] = ~(t[138] & t[139]);
  assign t[80] = ~(t[140]);
  assign t[81] = ~(t[141] & t[106]);
  assign t[82] = ~(x[7] & t[52]);
  assign t[83] = ~(t[141]);
  assign t[84] = ~(t[80]);
  assign t[85] = t[138] ? t[108] : t[107];
  assign t[86] = t[138] ? t[110] : t[109];
  assign t[87] = t[138] ? t[111] : t[81];
  assign t[88] = t[138] ? t[109] : t[110];
  assign t[89] = ~(t[157]);
  assign t[8] = ~(t[140] & t[141]);
  assign t[90] = ~(t[149] | t[150]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[112] & t[113]);
  assign t[93] = ~(t[158]);
  assign t[94] = ~(t[151] | t[152]);
  assign t[95] = ~(t[159]);
  assign t[96] = ~(t[160]);
  assign t[97] = ~(t[114] | t[115]);
  assign t[98] = ~(t[54] | t[116]);
  assign t[99] = ~(t[117] | t[118]);
  assign t[9] = ~(t[10] ^ t[12]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [163:0] x;
 output y;

 wire [635:0] t;
  assign t[0] = t[1] ? t[2] : t[388];
  assign t[100] = ~(t[411]);
  assign t[101] = ~(t[400] | t[401]);
  assign t[102] = ~(t[138] & t[140]);
  assign t[103] = ~(t[412]);
  assign t[104] = ~(t[413]);
  assign t[105] = ~(t[141] | t[142]);
  assign t[106] = ~(t[143] | t[144]);
  assign t[107] = ~(t[414] | t[145]);
  assign t[108] = t[391] ? x[94] : x[93];
  assign t[109] = ~(t[146] & t[147]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[415]);
  assign t[111] = ~(t[416]);
  assign t[112] = ~(t[148] | t[149]);
  assign t[113] = ~(t[150] | t[151]);
  assign t[114] = ~(t[417] | t[152]);
  assign t[115] = t[391] ? x[104] : x[103];
  assign t[116] = ~(t[146] & t[153]);
  assign t[117] = ~(t[122] | t[389]);
  assign t[118] = ~(t[154] & t[155]);
  assign t[119] = ~(t[390] | t[156]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = t[80] & t[389];
  assign t[121] = ~(t[122] | t[157]);
  assign t[122] = ~(t[391]);
  assign t[123] = t[389] ? t[159] : t[158];
  assign t[124] = ~(t[160] & t[392]);
  assign t[125] = ~(t[161] & t[156]);
  assign t[126] = ~(t[418]);
  assign t[127] = ~(t[405] | t[406]);
  assign t[128] = ~(t[162] & t[163]);
  assign t[129] = ~(t[164] & t[79]);
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = ~(t[80] | t[165]);
  assign t[131] = ~(t[80] | t[166]);
  assign t[132] = ~(t[419]);
  assign t[133] = ~(t[407] | t[408]);
  assign t[134] = ~(t[130] | t[167]);
  assign t[135] = ~(t[168] | t[169]);
  assign t[136] = ~(t[420]);
  assign t[137] = ~(t[409] | t[410]);
  assign t[138] = ~(t[49] | t[170]);
  assign t[139] = ~(t[171] | t[172]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = ~(t[167] | t[131]);
  assign t[141] = ~(t[421]);
  assign t[142] = ~(t[412] | t[413]);
  assign t[143] = ~(t[422]);
  assign t[144] = ~(t[423]);
  assign t[145] = ~(t[173] | t[174]);
  assign t[146] = ~(t[49] | t[175]);
  assign t[147] = ~(t[121] | t[176]);
  assign t[148] = ~(t[424]);
  assign t[149] = ~(t[415] | t[416]);
  assign t[14] = x[7] ? t[21] : t[20];
  assign t[150] = ~(t[425]);
  assign t[151] = ~(t[426]);
  assign t[152] = ~(t[177] | t[178]);
  assign t[153] = ~(t[179] | t[131]);
  assign t[154] = ~(t[392] & t[180]);
  assign t[155] = ~(x[7] & t[119]);
  assign t[156] = ~(t[392]);
  assign t[157] = t[389] ? t[158] : t[159];
  assign t[158] = ~(t[180] & t[156]);
  assign t[159] = ~(x[7] & t[181]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = x[7] & t[390];
  assign t[161] = ~(x[7] | t[390]);
  assign t[162] = ~(t[171] | t[182]);
  assign t[163] = ~(t[122] & t[183]);
  assign t[164] = ~(t[184] & t[185]);
  assign t[165] = t[389] ? t[124] : t[125];
  assign t[166] = t[389] ? t[187] : t[186];
  assign t[167] = ~(t[80] | t[188]);
  assign t[168] = t[172] | t[189];
  assign t[169] = ~(t[190] & t[79]);
  assign t[16] = x[7] ? t[25] : t[24];
  assign t[170] = ~(t[80] | t[191]);
  assign t[171] = ~(t[122] | t[192]);
  assign t[172] = ~(t[193] & t[77]);
  assign t[173] = ~(t[427]);
  assign t[174] = ~(t[422] | t[423]);
  assign t[175] = ~(t[134] & t[164]);
  assign t[176] = t[170] | t[194];
  assign t[177] = ~(t[428]);
  assign t[178] = ~(t[425] | t[426]);
  assign t[179] = ~(t[80] | t[195]);
  assign t[17] = ~(t[26] ^ t[27]);
  assign t[180] = ~(x[7] | t[196]);
  assign t[181] = ~(t[390] | t[392]);
  assign t[182] = ~(t[80] | t[197]);
  assign t[183] = ~(t[159] & t[154]);
  assign t[184] = t[392] & t[117];
  assign t[185] = t[161] | t[160];
  assign t[186] = ~(t[161] & t[392]);
  assign t[187] = ~(t[160] & t[156]);
  assign t[188] = t[389] ? t[159] : t[154];
  assign t[189] = ~(t[80] | t[198]);
  assign t[18] = t[28] ? x[21] : x[22];
  assign t[190] = ~(t[194] | t[179]);
  assign t[191] = t[389] ? t[186] : t[187];
  assign t[192] = t[389] ? t[125] : t[187];
  assign t[193] = ~(t[199] | t[121]);
  assign t[194] = ~(t[76]);
  assign t[195] = t[389] ? t[155] : t[158];
  assign t[196] = ~(t[390]);
  assign t[197] = t[389] ? t[158] : t[155];
  assign t[198] = t[389] ? t[154] : t[159];
  assign t[199] = ~(t[122] | t[200]);
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[389] ? t[187] : t[125];
  assign t[201] = t[1] ? t[202] : t[429];
  assign t[202] = x[6] ? t[204] : t[203];
  assign t[203] = x[7] ? t[206] : t[205];
  assign t[204] = t[207] ^ x[117];
  assign t[205] = t[208] ^ t[209];
  assign t[206] = ~(t[210] ^ t[211]);
  assign t[207] = x[118] ^ x[119];
  assign t[208] = t[391] ? x[118] : x[119];
  assign t[209] = ~(t[212] ^ t[213]);
  assign t[20] = ~(t[31] | t[32]);
  assign t[210] = x[7] ? t[215] : t[214];
  assign t[211] = ~(t[216] ^ t[217]);
  assign t[212] = x[7] ? t[219] : t[218];
  assign t[213] = ~(t[220] ^ t[221]);
  assign t[214] = ~(t[222] & t[223]);
  assign t[215] = t[224] ^ t[225];
  assign t[216] = x[7] ? t[227] : t[226];
  assign t[217] = x[7] ? t[229] : t[228];
  assign t[218] = ~(t[230] & t[231]);
  assign t[219] = t[232] ^ t[218];
  assign t[21] = ~(t[33] ^ t[34]);
  assign t[220] = x[7] ? t[234] : t[233];
  assign t[221] = x[7] ? t[236] : t[235];
  assign t[222] = ~(t[395] & t[51]);
  assign t[223] = ~(t[404] & t[237]);
  assign t[224] = t[238] ? x[121] : x[120];
  assign t[225] = ~(t[239] & t[240]);
  assign t[226] = ~(t[241] & t[242]);
  assign t[227] = t[243] ^ t[228];
  assign t[228] = ~(t[244] & t[245]);
  assign t[229] = t[246] ^ t[233];
  assign t[22] = x[7] ? t[36] : t[35];
  assign t[230] = ~(t[400] & t[64]);
  assign t[231] = ~(t[411] & t[247]);
  assign t[232] = t[391] ? x[123] : x[122];
  assign t[233] = ~(t[248] & t[249]);
  assign t[234] = t[250] ^ t[251];
  assign t[235] = ~(t[252] & t[253]);
  assign t[236] = t[254] ^ t[255];
  assign t[237] = ~(t[396] & t[50]);
  assign t[238] = ~(t[46]);
  assign t[239] = ~(t[405] & t[85]);
  assign t[23] = x[7] ? t[38] : t[37];
  assign t[240] = ~(t[418] & t[256]);
  assign t[241] = ~(t[409] & t[96]);
  assign t[242] = ~(t[420] & t[257]);
  assign t[243] = t[28] ? x[125] : x[124];
  assign t[244] = ~(t[407] & t[91]);
  assign t[245] = ~(t[419] & t[258]);
  assign t[246] = t[87] ? x[127] : x[126];
  assign t[247] = ~(t[401] & t[63]);
  assign t[248] = ~(t[415] & t[111]);
  assign t[249] = ~(t[424] & t[259]);
  assign t[24] = ~(t[39] | t[40]);
  assign t[250] = t[391] ? x[129] : x[128];
  assign t[251] = ~(t[260] & t[261]);
  assign t[252] = ~(t[412] & t[104]);
  assign t[253] = ~(t[421] & t[262]);
  assign t[254] = t[238] ? x[131] : x[130];
  assign t[255] = ~(t[263] & t[264]);
  assign t[256] = ~(t[406] & t[84]);
  assign t[257] = ~(t[410] & t[95]);
  assign t[258] = ~(t[408] & t[90]);
  assign t[259] = ~(t[416] & t[110]);
  assign t[25] = ~(t[24] ^ t[41]);
  assign t[260] = ~(t[425] & t[151]);
  assign t[261] = ~(t[428] & t[265]);
  assign t[262] = ~(t[413] & t[103]);
  assign t[263] = ~(t[422] & t[144]);
  assign t[264] = ~(t[427] & t[266]);
  assign t[265] = ~(t[426] & t[150]);
  assign t[266] = ~(t[423] & t[143]);
  assign t[267] = t[1] ? t[268] : t[430];
  assign t[268] = x[6] ? t[270] : t[269];
  assign t[269] = x[7] ? t[272] : t[271];
  assign t[26] = x[7] ? t[43] : t[42];
  assign t[270] = t[273] ^ x[133];
  assign t[271] = t[274] ^ t[275];
  assign t[272] = ~(t[276] ^ t[277]);
  assign t[273] = x[134] ^ x[135];
  assign t[274] = t[391] ? x[134] : x[135];
  assign t[275] = ~(t[278] ^ t[279]);
  assign t[276] = x[7] ? t[281] : t[280];
  assign t[277] = ~(t[282] ^ t[283]);
  assign t[278] = x[7] ? t[285] : t[284];
  assign t[279] = ~(t[286] ^ t[287]);
  assign t[27] = x[7] ? t[45] : t[44];
  assign t[280] = ~(t[288] & t[289]);
  assign t[281] = t[290] ^ t[291];
  assign t[282] = x[7] ? t[293] : t[292];
  assign t[283] = x[7] ? t[295] : t[294];
  assign t[284] = ~(t[296] & t[297]);
  assign t[285] = t[298] ^ t[284];
  assign t[286] = x[7] ? t[300] : t[299];
  assign t[287] = x[7] ? t[302] : t[301];
  assign t[288] = ~(t[51] & t[82]);
  assign t[289] = ~(t[303] & t[393]);
  assign t[28] = ~(t[46]);
  assign t[290] = t[87] ? x[137] : x[136];
  assign t[291] = ~(t[304] & t[305]);
  assign t[292] = ~(t[306] & t[307]);
  assign t[293] = t[308] ^ t[299];
  assign t[294] = ~(t[309] & t[310]);
  assign t[295] = t[311] ^ t[292];
  assign t[296] = ~(t[64] & t[100]);
  assign t[297] = ~(t[312] & t[394]);
  assign t[298] = t[391] ? x[139] : x[138];
  assign t[299] = ~(t[313] & t[314]);
  assign t[29] = ~(t[47] | t[48]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = t[315] ^ t[316];
  assign t[301] = ~(t[317] & t[318]);
  assign t[302] = t[319] ^ t[320];
  assign t[303] = ~(t[321] & t[50]);
  assign t[304] = ~(t[85] & t[126]);
  assign t[305] = ~(t[322] & t[397]);
  assign t[306] = ~(t[91] & t[132]);
  assign t[307] = ~(t[323] & t[398]);
  assign t[308] = t[87] ? x[141] : x[140];
  assign t[309] = ~(t[96] & t[136]);
  assign t[30] = ~(t[49]);
  assign t[310] = ~(t[324] & t[399]);
  assign t[311] = t[391] ? x[143] : x[142];
  assign t[312] = ~(t[325] & t[63]);
  assign t[313] = ~(t[111] & t[148]);
  assign t[314] = ~(t[326] & t[403]);
  assign t[315] = t[391] ? x[145] : x[144];
  assign t[316] = ~(t[327] & t[328]);
  assign t[317] = ~(t[104] & t[141]);
  assign t[318] = ~(t[329] & t[402]);
  assign t[319] = t[87] ? x[147] : x[146];
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = ~(t[330] & t[331]);
  assign t[321] = ~(t[404] & t[396]);
  assign t[322] = ~(t[332] & t[84]);
  assign t[323] = ~(t[333] & t[90]);
  assign t[324] = ~(t[334] & t[95]);
  assign t[325] = ~(t[411] & t[401]);
  assign t[326] = ~(t[335] & t[110]);
  assign t[327] = ~(t[151] & t[177]);
  assign t[328] = ~(t[336] & t[417]);
  assign t[329] = ~(t[337] & t[103]);
  assign t[32] = ~(t[393] | t[52]);
  assign t[330] = ~(t[144] & t[173]);
  assign t[331] = ~(t[338] & t[414]);
  assign t[332] = ~(t[418] & t[406]);
  assign t[333] = ~(t[419] & t[408]);
  assign t[334] = ~(t[420] & t[410]);
  assign t[335] = ~(t[424] & t[416]);
  assign t[336] = ~(t[339] & t[150]);
  assign t[337] = ~(t[421] & t[413]);
  assign t[338] = ~(t[340] & t[143]);
  assign t[339] = ~(t[428] & t[426]);
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = ~(t[427] & t[423]);
  assign t[341] = t[1] ? t[342] : t[431];
  assign t[342] = x[6] ? t[344] : t[343];
  assign t[343] = x[7] ? t[346] : t[345];
  assign t[344] = t[347] ^ x[149];
  assign t[345] = t[348] ^ t[349];
  assign t[346] = ~(t[350] ^ t[351]);
  assign t[347] = x[150] ^ x[151];
  assign t[348] = t[391] ? x[150] : x[151];
  assign t[349] = ~(t[352] ^ t[353]);
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[350] = x[7] ? t[355] : t[354];
  assign t[351] = ~(t[356] ^ t[357]);
  assign t[352] = x[7] ? t[359] : t[358];
  assign t[353] = ~(t[360] ^ t[361]);
  assign t[354] = ~(t[288] & t[362]);
  assign t[355] = t[363] ^ t[364];
  assign t[356] = x[7] ? t[366] : t[365];
  assign t[357] = x[7] ? t[368] : t[367];
  assign t[358] = ~(t[296] & t[369]);
  assign t[359] = t[370] ^ t[358];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = x[7] ? t[372] : t[371];
  assign t[361] = x[7] ? t[374] : t[373];
  assign t[362] = t[31] | t[393];
  assign t[363] = t[87] ? x[153] : x[152];
  assign t[364] = ~(t[304] & t[375]);
  assign t[365] = ~(t[306] & t[376]);
  assign t[366] = t[377] ^ t[371];
  assign t[367] = ~(t[309] & t[378]);
  assign t[368] = t[379] ^ t[365];
  assign t[369] = t[39] | t[394];
  assign t[36] = ~(t[44] ^ t[59]);
  assign t[370] = t[391] ? x[155] : x[154];
  assign t[371] = ~(t[313] & t[380]);
  assign t[372] = t[381] ^ t[382];
  assign t[373] = ~(t[317] & t[383]);
  assign t[374] = t[384] ^ t[385];
  assign t[375] = t[53] | t[397];
  assign t[376] = t[57] | t[398];
  assign t[377] = t[87] ? x[157] : x[156];
  assign t[378] = t[60] | t[399];
  assign t[379] = t[87] ? x[159] : x[158];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[72] | t[403];
  assign t[381] = t[391] ? x[161] : x[160];
  assign t[382] = ~(t[327] & t[386]);
  assign t[383] = t[68] | t[402];
  assign t[384] = t[28] ? x[163] : x[162];
  assign t[385] = ~(t[330] & t[387]);
  assign t[386] = t[113] | t[417];
  assign t[387] = t[106] | t[414];
  assign t[388] = (t[432]);
  assign t[389] = (t[433]);
  assign t[38] = ~(t[35] ^ t[62]);
  assign t[390] = (t[434]);
  assign t[391] = (t[435]);
  assign t[392] = (t[436]);
  assign t[393] = (t[437]);
  assign t[394] = (t[438]);
  assign t[395] = (t[439]);
  assign t[396] = (t[440]);
  assign t[397] = (t[441]);
  assign t[398] = (t[442]);
  assign t[399] = (t[443]);
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (t[444]);
  assign t[401] = (t[445]);
  assign t[402] = (t[446]);
  assign t[403] = (t[447]);
  assign t[404] = (t[448]);
  assign t[405] = (t[449]);
  assign t[406] = (t[450]);
  assign t[407] = (t[451]);
  assign t[408] = (t[452]);
  assign t[409] = (t[453]);
  assign t[40] = ~(t[394] | t[65]);
  assign t[410] = (t[454]);
  assign t[411] = (t[455]);
  assign t[412] = (t[456]);
  assign t[413] = (t[457]);
  assign t[414] = (t[458]);
  assign t[415] = (t[459]);
  assign t[416] = (t[460]);
  assign t[417] = (t[461]);
  assign t[418] = (t[462]);
  assign t[419] = (t[463]);
  assign t[41] = ~(t[66] ^ t[67]);
  assign t[420] = (t[464]);
  assign t[421] = (t[465]);
  assign t[422] = (t[466]);
  assign t[423] = (t[467]);
  assign t[424] = (t[468]);
  assign t[425] = (t[469]);
  assign t[426] = (t[470]);
  assign t[427] = (t[471]);
  assign t[428] = (t[472]);
  assign t[429] = (t[473]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (t[474]);
  assign t[431] = (t[475]);
  assign t[432] = t[476] ^ x[5];
  assign t[433] = t[477] ^ x[11];
  assign t[434] = t[478] ^ x[14];
  assign t[435] = t[479] ^ x[17];
  assign t[436] = t[480] ^ x[20];
  assign t[437] = t[481] ^ x[28];
  assign t[438] = t[482] ^ x[34];
  assign t[439] = t[483] ^ x[35];
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = t[484] ^ x[36];
  assign t[441] = t[485] ^ x[42];
  assign t[442] = t[486] ^ x[50];
  assign t[443] = t[487] ^ x[56];
  assign t[444] = t[488] ^ x[57];
  assign t[445] = t[489] ^ x[58];
  assign t[446] = t[490] ^ x[66];
  assign t[447] = t[491] ^ x[72];
  assign t[448] = t[492] ^ x[73];
  assign t[449] = t[493] ^ x[74];
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = t[494] ^ x[75];
  assign t[451] = t[495] ^ x[76];
  assign t[452] = t[496] ^ x[77];
  assign t[453] = t[497] ^ x[80];
  assign t[454] = t[498] ^ x[81];
  assign t[455] = t[499] ^ x[84];
  assign t[456] = t[500] ^ x[85];
  assign t[457] = t[501] ^ x[86];
  assign t[458] = t[502] ^ x[92];
  assign t[459] = t[503] ^ x[95];
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[460] = t[504] ^ x[96];
  assign t[461] = t[505] ^ x[102];
  assign t[462] = t[506] ^ x[105];
  assign t[463] = t[507] ^ x[106];
  assign t[464] = t[508] ^ x[107];
  assign t[465] = t[509] ^ x[108];
  assign t[466] = t[510] ^ x[109];
  assign t[467] = t[511] ^ x[110];
  assign t[468] = t[512] ^ x[111];
  assign t[469] = t[513] ^ x[112];
  assign t[46] = ~(t[391]);
  assign t[470] = t[514] ^ x[113];
  assign t[471] = t[515] ^ x[114];
  assign t[472] = t[516] ^ x[115];
  assign t[473] = t[517] ^ x[116];
  assign t[474] = t[518] ^ x[132];
  assign t[475] = t[519] ^ x[148];
  assign t[476] = (~t[520] & t[521]);
  assign t[477] = (~t[522] & t[523]);
  assign t[478] = (~t[524] & t[525]);
  assign t[479] = (~t[526] & t[527]);
  assign t[47] = ~(t[76] & t[77]);
  assign t[480] = (~t[528] & t[529]);
  assign t[481] = (~t[530] & t[531]);
  assign t[482] = (~t[532] & t[533]);
  assign t[483] = (~t[530] & t[534]);
  assign t[484] = (~t[530] & t[535]);
  assign t[485] = (~t[536] & t[537]);
  assign t[486] = (~t[538] & t[539]);
  assign t[487] = (~t[540] & t[541]);
  assign t[488] = (~t[532] & t[542]);
  assign t[489] = (~t[532] & t[543]);
  assign t[48] = ~(t[78] & t[79]);
  assign t[490] = (~t[544] & t[545]);
  assign t[491] = (~t[546] & t[547]);
  assign t[492] = (~t[530] & t[548]);
  assign t[493] = (~t[536] & t[549]);
  assign t[494] = (~t[536] & t[550]);
  assign t[495] = (~t[538] & t[551]);
  assign t[496] = (~t[538] & t[552]);
  assign t[497] = (~t[540] & t[553]);
  assign t[498] = (~t[540] & t[554]);
  assign t[499] = (~t[532] & t[555]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = ~(x[6]);
  assign t[500] = (~t[544] & t[556]);
  assign t[501] = (~t[544] & t[557]);
  assign t[502] = (~t[558] & t[559]);
  assign t[503] = (~t[546] & t[560]);
  assign t[504] = (~t[546] & t[561]);
  assign t[505] = (~t[562] & t[563]);
  assign t[506] = (~t[536] & t[564]);
  assign t[507] = (~t[538] & t[565]);
  assign t[508] = (~t[540] & t[566]);
  assign t[509] = (~t[544] & t[567]);
  assign t[50] = ~(t[395]);
  assign t[510] = (~t[558] & t[568]);
  assign t[511] = (~t[558] & t[569]);
  assign t[512] = (~t[546] & t[570]);
  assign t[513] = (~t[562] & t[571]);
  assign t[514] = (~t[562] & t[572]);
  assign t[515] = (~t[558] & t[573]);
  assign t[516] = (~t[562] & t[574]);
  assign t[517] = (~t[520] & t[575]);
  assign t[518] = (~t[520] & t[576]);
  assign t[519] = (~t[520] & t[577]);
  assign t[51] = ~(t[396]);
  assign t[520] = t[578] ^ x[4];
  assign t[521] = t[579] ^ x[5];
  assign t[522] = t[580] ^ x[10];
  assign t[523] = t[581] ^ x[11];
  assign t[524] = t[582] ^ x[13];
  assign t[525] = t[583] ^ x[14];
  assign t[526] = t[584] ^ x[16];
  assign t[527] = t[585] ^ x[17];
  assign t[528] = t[586] ^ x[19];
  assign t[529] = t[587] ^ x[20];
  assign t[52] = ~(t[82] | t[83]);
  assign t[530] = t[588] ^ x[27];
  assign t[531] = t[589] ^ x[28];
  assign t[532] = t[590] ^ x[33];
  assign t[533] = t[591] ^ x[34];
  assign t[534] = t[592] ^ x[35];
  assign t[535] = t[593] ^ x[36];
  assign t[536] = t[594] ^ x[41];
  assign t[537] = t[595] ^ x[42];
  assign t[538] = t[596] ^ x[49];
  assign t[539] = t[597] ^ x[50];
  assign t[53] = ~(t[84] | t[85]);
  assign t[540] = t[598] ^ x[55];
  assign t[541] = t[599] ^ x[56];
  assign t[542] = t[600] ^ x[57];
  assign t[543] = t[601] ^ x[58];
  assign t[544] = t[602] ^ x[65];
  assign t[545] = t[603] ^ x[66];
  assign t[546] = t[604] ^ x[71];
  assign t[547] = t[605] ^ x[72];
  assign t[548] = t[606] ^ x[73];
  assign t[549] = t[607] ^ x[74];
  assign t[54] = ~(t[397] | t[86]);
  assign t[550] = t[608] ^ x[75];
  assign t[551] = t[609] ^ x[76];
  assign t[552] = t[610] ^ x[77];
  assign t[553] = t[611] ^ x[80];
  assign t[554] = t[612] ^ x[81];
  assign t[555] = t[613] ^ x[84];
  assign t[556] = t[614] ^ x[85];
  assign t[557] = t[615] ^ x[86];
  assign t[558] = t[616] ^ x[91];
  assign t[559] = t[617] ^ x[92];
  assign t[55] = t[87] ? x[44] : x[43];
  assign t[560] = t[618] ^ x[95];
  assign t[561] = t[619] ^ x[96];
  assign t[562] = t[620] ^ x[101];
  assign t[563] = t[621] ^ x[102];
  assign t[564] = t[622] ^ x[105];
  assign t[565] = t[623] ^ x[106];
  assign t[566] = t[624] ^ x[107];
  assign t[567] = t[625] ^ x[108];
  assign t[568] = t[626] ^ x[109];
  assign t[569] = t[627] ^ x[110];
  assign t[56] = ~(t[88] & t[89]);
  assign t[570] = t[628] ^ x[111];
  assign t[571] = t[629] ^ x[112];
  assign t[572] = t[630] ^ x[113];
  assign t[573] = t[631] ^ x[114];
  assign t[574] = t[632] ^ x[115];
  assign t[575] = t[633] ^ x[116];
  assign t[576] = t[634] ^ x[132];
  assign t[577] = t[635] ^ x[148];
  assign t[578] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[579] = (x[0]);
  assign t[57] = ~(t[90] | t[91]);
  assign t[580] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[581] = (x[9]);
  assign t[582] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[583] = (x[12]);
  assign t[584] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[585] = (x[15]);
  assign t[586] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[587] = (x[18]);
  assign t[588] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[589] = (x[24]);
  assign t[58] = ~(t[398] | t[92]);
  assign t[590] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[591] = (x[30]);
  assign t[592] = (x[25]);
  assign t[593] = (x[26]);
  assign t[594] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[595] = (x[38]);
  assign t[596] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[597] = (x[46]);
  assign t[598] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[599] = (x[52]);
  assign t[59] = ~(t[93] ^ t[94]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[600] = (x[31]);
  assign t[601] = (x[32]);
  assign t[602] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[603] = (x[62]);
  assign t[604] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[605] = (x[68]);
  assign t[606] = (x[23]);
  assign t[607] = (x[39]);
  assign t[608] = (x[40]);
  assign t[609] = (x[47]);
  assign t[60] = ~(t[95] | t[96]);
  assign t[610] = (x[48]);
  assign t[611] = (x[53]);
  assign t[612] = (x[54]);
  assign t[613] = (x[29]);
  assign t[614] = (x[63]);
  assign t[615] = (x[64]);
  assign t[616] = (x[87] & ~x[88] & ~x[89] & ~x[90]) | (~x[87] & x[88] & ~x[89] & ~x[90]) | (~x[87] & ~x[88] & x[89] & ~x[90]) | (~x[87] & ~x[88] & ~x[89] & x[90]) | (x[87] & x[88] & x[89] & ~x[90]) | (x[87] & x[88] & ~x[89] & x[90]) | (x[87] & ~x[88] & x[89] & x[90]) | (~x[87] & x[88] & x[89] & x[90]);
  assign t[617] = (x[88]);
  assign t[618] = (x[69]);
  assign t[619] = (x[70]);
  assign t[61] = ~(t[399] | t[97]);
  assign t[620] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[621] = (x[98]);
  assign t[622] = (x[37]);
  assign t[623] = (x[45]);
  assign t[624] = (x[51]);
  assign t[625] = (x[61]);
  assign t[626] = (x[89]);
  assign t[627] = (x[90]);
  assign t[628] = (x[67]);
  assign t[629] = (x[99]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[630] = (x[100]);
  assign t[631] = (x[87]);
  assign t[632] = (x[97]);
  assign t[633] = (x[1]);
  assign t[634] = (x[2]);
  assign t[635] = (x[3]);
  assign t[63] = ~(t[400]);
  assign t[64] = ~(t[401]);
  assign t[65] = ~(t[100] | t[101]);
  assign t[66] = t[391] ? x[60] : x[59];
  assign t[67] = t[47] | t[102];
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = ~(t[402] | t[105]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[108] ^ t[109]);
  assign t[72] = ~(t[110] | t[111]);
  assign t[73] = ~(t[403] | t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[115] ^ t[116]);
  assign t[76] = ~(t[117] & t[118]);
  assign t[77] = ~(t[119] & t[120]);
  assign t[78] = ~(t[121]);
  assign t[79] = t[122] | t[123];
  assign t[7] = ~(t[389] & t[390]);
  assign t[80] = ~(t[122]);
  assign t[81] = t[389] ? t[125] : t[124];
  assign t[82] = ~(t[404]);
  assign t[83] = ~(t[395] | t[396]);
  assign t[84] = ~(t[405]);
  assign t[85] = ~(t[406]);
  assign t[86] = ~(t[126] | t[127]);
  assign t[87] = ~(t[46]);
  assign t[88] = ~(t[128] | t[129]);
  assign t[89] = ~(t[130] | t[131]);
  assign t[8] = ~(t[391] & t[392]);
  assign t[90] = ~(t[407]);
  assign t[91] = ~(t[408]);
  assign t[92] = ~(t[132] | t[133]);
  assign t[93] = t[87] ? x[79] : x[78];
  assign t[94] = ~(t[134] & t[135]);
  assign t[95] = ~(t[409]);
  assign t[96] = ~(t[410]);
  assign t[97] = ~(t[136] | t[137]);
  assign t[98] = t[87] ? x[83] : x[82];
  assign t[99] = ~(t[138] & t[139]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0] & ~t[201] & ~t[267] & ~t[341]) | (~t[0] & t[201] & ~t[267] & ~t[341]) | (~t[0] & ~t[201] & t[267] & ~t[341]) | (~t[0] & ~t[201] & ~t[267] & t[341]) | (t[0] & t[201] & t[267] & ~t[341]) | (t[0] & t[201] & ~t[267] & t[341]) | (t[0] & ~t[201] & t[267] & t[341]) | (~t[0] & t[201] & t[267] & t[341]);
endmodule

module R2ind126(x, y);
 input [115:0] x;
 output y;

 wire [332:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[141]);
  assign t[101] = (t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[103] ? x[21] : x[22];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = t[182] ^ x[5];
  assign t[142] = t[183] ^ x[11];
  assign t[143] = t[184] ^ x[14];
  assign t[144] = t[185] ^ x[17];
  assign t[145] = t[186] ^ x[20];
  assign t[146] = t[187] ^ x[28];
  assign t[147] = t[188] ^ x[36];
  assign t[148] = t[189] ^ x[39];
  assign t[149] = t[190] ^ x[40];
  assign t[14] = x[7] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[46];
  assign t[151] = t[192] ^ x[52];
  assign t[152] = t[193] ^ x[60];
  assign t[153] = t[194] ^ x[63];
  assign t[154] = t[195] ^ x[64];
  assign t[155] = t[196] ^ x[70];
  assign t[156] = t[197] ^ x[78];
  assign t[157] = t[198] ^ x[81];
  assign t[158] = t[199] ^ x[82];
  assign t[159] = t[200] ^ x[83];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[84];
  assign t[161] = t[202] ^ x[85];
  assign t[162] = t[203] ^ x[86];
  assign t[163] = t[204] ^ x[87];
  assign t[164] = t[205] ^ x[88];
  assign t[165] = t[206] ^ x[89];
  assign t[166] = t[207] ^ x[90];
  assign t[167] = t[208] ^ x[96];
  assign t[168] = t[209] ^ x[97];
  assign t[169] = t[210] ^ x[98];
  assign t[16] = x[7] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[104];
  assign t[171] = t[212] ^ x[105];
  assign t[172] = t[213] ^ x[106];
  assign t[173] = t[214] ^ x[107];
  assign t[174] = t[215] ^ x[108];
  assign t[175] = t[216] ^ x[109];
  assign t[176] = t[217] ^ x[110];
  assign t[177] = t[218] ^ x[111];
  assign t[178] = t[219] ^ x[112];
  assign t[179] = t[220] ^ x[113];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[114];
  assign t[181] = t[222] ^ x[115];
  assign t[182] = (~t[223] & t[224]);
  assign t[183] = (~t[225] & t[226]);
  assign t[184] = (~t[227] & t[228]);
  assign t[185] = (~t[229] & t[230]);
  assign t[186] = (~t[231] & t[232]);
  assign t[187] = (~t[233] & t[234]);
  assign t[188] = (~t[235] & t[236]);
  assign t[189] = (~t[233] & t[237]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (~t[233] & t[238]);
  assign t[191] = (~t[239] & t[240]);
  assign t[192] = (~t[241] & t[242]);
  assign t[193] = (~t[243] & t[244]);
  assign t[194] = (~t[235] & t[245]);
  assign t[195] = (~t[235] & t[246]);
  assign t[196] = (~t[247] & t[248]);
  assign t[197] = (~t[249] & t[250]);
  assign t[198] = (~t[233] & t[251]);
  assign t[199] = (~t[239] & t[252]);
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (~t[239] & t[253]);
  assign t[201] = (~t[241] & t[254]);
  assign t[202] = (~t[241] & t[255]);
  assign t[203] = (~t[243] & t[256]);
  assign t[204] = (~t[243] & t[257]);
  assign t[205] = (~t[235] & t[258]);
  assign t[206] = (~t[247] & t[259]);
  assign t[207] = (~t[247] & t[260]);
  assign t[208] = (~t[261] & t[262]);
  assign t[209] = (~t[249] & t[263]);
  assign t[20] = x[7] ? t[31] : t[30];
  assign t[210] = (~t[249] & t[264]);
  assign t[211] = (~t[265] & t[266]);
  assign t[212] = (~t[239] & t[267]);
  assign t[213] = (~t[241] & t[268]);
  assign t[214] = (~t[243] & t[269]);
  assign t[215] = (~t[247] & t[270]);
  assign t[216] = (~t[261] & t[271]);
  assign t[217] = (~t[261] & t[272]);
  assign t[218] = (~t[249] & t[273]);
  assign t[219] = (~t[265] & t[274]);
  assign t[21] = x[7] ? t[33] : t[32];
  assign t[220] = (~t[265] & t[275]);
  assign t[221] = (~t[261] & t[276]);
  assign t[222] = (~t[265] & t[277]);
  assign t[223] = t[278] ^ x[4];
  assign t[224] = t[279] ^ x[5];
  assign t[225] = t[280] ^ x[10];
  assign t[226] = t[281] ^ x[11];
  assign t[227] = t[282] ^ x[13];
  assign t[228] = t[283] ^ x[14];
  assign t[229] = t[284] ^ x[16];
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = t[285] ^ x[17];
  assign t[231] = t[286] ^ x[19];
  assign t[232] = t[287] ^ x[20];
  assign t[233] = t[288] ^ x[27];
  assign t[234] = t[289] ^ x[28];
  assign t[235] = t[290] ^ x[35];
  assign t[236] = t[291] ^ x[36];
  assign t[237] = t[292] ^ x[39];
  assign t[238] = t[293] ^ x[40];
  assign t[239] = t[294] ^ x[45];
  assign t[23] = t[36] ^ t[22];
  assign t[240] = t[295] ^ x[46];
  assign t[241] = t[296] ^ x[51];
  assign t[242] = t[297] ^ x[52];
  assign t[243] = t[298] ^ x[59];
  assign t[244] = t[299] ^ x[60];
  assign t[245] = t[300] ^ x[63];
  assign t[246] = t[301] ^ x[64];
  assign t[247] = t[302] ^ x[69];
  assign t[248] = t[303] ^ x[70];
  assign t[249] = t[304] ^ x[77];
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = t[305] ^ x[78];
  assign t[251] = t[306] ^ x[81];
  assign t[252] = t[307] ^ x[82];
  assign t[253] = t[308] ^ x[83];
  assign t[254] = t[309] ^ x[84];
  assign t[255] = t[310] ^ x[85];
  assign t[256] = t[311] ^ x[86];
  assign t[257] = t[312] ^ x[87];
  assign t[258] = t[313] ^ x[88];
  assign t[259] = t[314] ^ x[89];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[315] ^ x[90];
  assign t[261] = t[316] ^ x[95];
  assign t[262] = t[317] ^ x[96];
  assign t[263] = t[318] ^ x[97];
  assign t[264] = t[319] ^ x[98];
  assign t[265] = t[320] ^ x[103];
  assign t[266] = t[321] ^ x[104];
  assign t[267] = t[322] ^ x[105];
  assign t[268] = t[323] ^ x[106];
  assign t[269] = t[324] ^ x[107];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[325] ^ x[108];
  assign t[271] = t[326] ^ x[109];
  assign t[272] = t[327] ^ x[110];
  assign t[273] = t[328] ^ x[111];
  assign t[274] = t[329] ^ x[112];
  assign t[275] = t[330] ^ x[113];
  assign t[276] = t[331] ^ x[114];
  assign t[277] = t[332] ^ x[115];
  assign t[278] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[279] = (x[3]);
  assign t[27] = t[43] | t[105];
  assign t[280] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[281] = (x[9]);
  assign t[282] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[283] = (x[12]);
  assign t[284] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[285] = (x[15]);
  assign t[286] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[287] = (x[18]);
  assign t[288] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[289] = (x[24]);
  assign t[28] = t[44] ? x[30] : x[29];
  assign t[290] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[291] = (x[32]);
  assign t[292] = (x[26]);
  assign t[293] = (x[23]);
  assign t[294] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[295] = (x[42]);
  assign t[296] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[297] = (x[48]);
  assign t[298] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[299] = (x[56]);
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = (x[34]);
  assign t[301] = (x[31]);
  assign t[302] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[303] = (x[66]);
  assign t[304] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[305] = (x[74]);
  assign t[306] = (x[25]);
  assign t[307] = (x[44]);
  assign t[308] = (x[41]);
  assign t[309] = (x[50]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[310] = (x[47]);
  assign t[311] = (x[58]);
  assign t[312] = (x[55]);
  assign t[313] = (x[33]);
  assign t[314] = (x[68]);
  assign t[315] = (x[65]);
  assign t[316] = (x[91] & ~x[92] & ~x[93] & ~x[94]) | (~x[91] & x[92] & ~x[93] & ~x[94]) | (~x[91] & ~x[92] & x[93] & ~x[94]) | (~x[91] & ~x[92] & ~x[93] & x[94]) | (x[91] & x[92] & x[93] & ~x[94]) | (x[91] & x[92] & ~x[93] & x[94]) | (x[91] & ~x[92] & x[93] & x[94]) | (~x[91] & x[92] & x[93] & x[94]);
  assign t[317] = (x[92]);
  assign t[318] = (x[76]);
  assign t[319] = (x[73]);
  assign t[31] = t[49] ^ t[37];
  assign t[320] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[321] = (x[100]);
  assign t[322] = (x[43]);
  assign t[323] = (x[49]);
  assign t[324] = (x[57]);
  assign t[325] = (x[67]);
  assign t[326] = (x[94]);
  assign t[327] = (x[91]);
  assign t[328] = (x[75]);
  assign t[329] = (x[102]);
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = (x[99]);
  assign t[331] = (x[93]);
  assign t[332] = (x[101]);
  assign t[33] = t[52] ^ t[30];
  assign t[34] = ~(t[53] & t[54]);
  assign t[35] = t[55] | t[106];
  assign t[36] = t[103] ? x[38] : x[37];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[107]);
  assign t[42] = ~(t[108]);
  assign t[43] = ~(t[64] | t[41]);
  assign t[44] = ~(t[65]);
  assign t[45] = ~(t[66] & t[67]);
  assign t[46] = t[68] | t[109];
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = t[71] | t[110];
  assign t[49] = t[44] ? x[54] : x[53];
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[111];
  assign t[52] = t[44] ? x[62] : x[61];
  assign t[53] = ~(t[112]);
  assign t[54] = ~(t[113]);
  assign t[55] = ~(t[75] | t[53]);
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = t[78] | t[114];
  assign t[58] = t[103] ? x[72] : x[71];
  assign t[59] = ~(t[79] & t[80]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[115];
  assign t[62] = t[84] ? x[80] : x[79];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = ~(t[116]);
  assign t[65] = ~(t[103]);
  assign t[66] = ~(t[117]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[87] | t[66]);
  assign t[69] = ~(t[119]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[120]);
  assign t[71] = ~(t[88] | t[69]);
  assign t[72] = ~(t[121]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[89] | t[72]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[90] | t[76]);
  assign t[79] = ~(t[91] & t[92]);
  assign t[7] = ~(t[101] & t[102]);
  assign t[80] = t[93] | t[126];
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[94] | t[81]);
  assign t[84] = ~(t[65]);
  assign t[85] = ~(t[95] & t[96]);
  assign t[86] = t[97] | t[129];
  assign t[87] = ~(t[130]);
  assign t[88] = ~(t[131]);
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[103] & t[104]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[98] | t[91]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[99] | t[95]);
  assign t[98] = ~(t[139]);
  assign t[99] = ~(t[140]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [115:0] x;
 output y;

 wire [340:0] t;
  assign t[0] = t[1] ? t[2] : t[108];
  assign t[100] = ~(t[144]);
  assign t[101] = ~(t[145]);
  assign t[102] = ~(t[146]);
  assign t[103] = ~(t[106] & t[107]);
  assign t[104] = ~(t[143] & t[142]);
  assign t[105] = ~(t[147]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[111] ? x[21] : x[22];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = t[190] ^ x[5];
  assign t[14] = x[7] ? t[19] : t[18];
  assign t[150] = t[191] ^ x[11];
  assign t[151] = t[192] ^ x[14];
  assign t[152] = t[193] ^ x[17];
  assign t[153] = t[194] ^ x[20];
  assign t[154] = t[195] ^ x[28];
  assign t[155] = t[196] ^ x[36];
  assign t[156] = t[197] ^ x[39];
  assign t[157] = t[198] ^ x[40];
  assign t[158] = t[199] ^ x[46];
  assign t[159] = t[200] ^ x[52];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[201] ^ x[60];
  assign t[161] = t[202] ^ x[63];
  assign t[162] = t[203] ^ x[64];
  assign t[163] = t[204] ^ x[70];
  assign t[164] = t[205] ^ x[78];
  assign t[165] = t[206] ^ x[81];
  assign t[166] = t[207] ^ x[82];
  assign t[167] = t[208] ^ x[83];
  assign t[168] = t[209] ^ x[84];
  assign t[169] = t[210] ^ x[85];
  assign t[16] = x[7] ? t[23] : t[22];
  assign t[170] = t[211] ^ x[86];
  assign t[171] = t[212] ^ x[87];
  assign t[172] = t[213] ^ x[88];
  assign t[173] = t[214] ^ x[89];
  assign t[174] = t[215] ^ x[90];
  assign t[175] = t[216] ^ x[96];
  assign t[176] = t[217] ^ x[97];
  assign t[177] = t[218] ^ x[98];
  assign t[178] = t[219] ^ x[104];
  assign t[179] = t[220] ^ x[105];
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = t[221] ^ x[106];
  assign t[181] = t[222] ^ x[107];
  assign t[182] = t[223] ^ x[108];
  assign t[183] = t[224] ^ x[109];
  assign t[184] = t[225] ^ x[110];
  assign t[185] = t[226] ^ x[111];
  assign t[186] = t[227] ^ x[112];
  assign t[187] = t[228] ^ x[113];
  assign t[188] = t[229] ^ x[114];
  assign t[189] = t[230] ^ x[115];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = (~t[231] & t[232]);
  assign t[191] = (~t[233] & t[234]);
  assign t[192] = (~t[235] & t[236]);
  assign t[193] = (~t[237] & t[238]);
  assign t[194] = (~t[239] & t[240]);
  assign t[195] = (~t[241] & t[242]);
  assign t[196] = (~t[243] & t[244]);
  assign t[197] = (~t[241] & t[245]);
  assign t[198] = (~t[241] & t[246]);
  assign t[199] = (~t[247] & t[248]);
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (~t[249] & t[250]);
  assign t[201] = (~t[251] & t[252]);
  assign t[202] = (~t[243] & t[253]);
  assign t[203] = (~t[243] & t[254]);
  assign t[204] = (~t[255] & t[256]);
  assign t[205] = (~t[257] & t[258]);
  assign t[206] = (~t[241] & t[259]);
  assign t[207] = (~t[247] & t[260]);
  assign t[208] = (~t[247] & t[261]);
  assign t[209] = (~t[249] & t[262]);
  assign t[20] = x[7] ? t[31] : t[30];
  assign t[210] = (~t[249] & t[263]);
  assign t[211] = (~t[251] & t[264]);
  assign t[212] = (~t[251] & t[265]);
  assign t[213] = (~t[243] & t[266]);
  assign t[214] = (~t[255] & t[267]);
  assign t[215] = (~t[255] & t[268]);
  assign t[216] = (~t[269] & t[270]);
  assign t[217] = (~t[257] & t[271]);
  assign t[218] = (~t[257] & t[272]);
  assign t[219] = (~t[273] & t[274]);
  assign t[21] = x[7] ? t[33] : t[32];
  assign t[220] = (~t[247] & t[275]);
  assign t[221] = (~t[249] & t[276]);
  assign t[222] = (~t[251] & t[277]);
  assign t[223] = (~t[255] & t[278]);
  assign t[224] = (~t[269] & t[279]);
  assign t[225] = (~t[269] & t[280]);
  assign t[226] = (~t[257] & t[281]);
  assign t[227] = (~t[273] & t[282]);
  assign t[228] = (~t[273] & t[283]);
  assign t[229] = (~t[269] & t[284]);
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = (~t[273] & t[285]);
  assign t[231] = t[286] ^ x[4];
  assign t[232] = t[287] ^ x[5];
  assign t[233] = t[288] ^ x[10];
  assign t[234] = t[289] ^ x[11];
  assign t[235] = t[290] ^ x[13];
  assign t[236] = t[291] ^ x[14];
  assign t[237] = t[292] ^ x[16];
  assign t[238] = t[293] ^ x[17];
  assign t[239] = t[294] ^ x[19];
  assign t[23] = t[36] ^ t[22];
  assign t[240] = t[295] ^ x[20];
  assign t[241] = t[296] ^ x[27];
  assign t[242] = t[297] ^ x[28];
  assign t[243] = t[298] ^ x[35];
  assign t[244] = t[299] ^ x[36];
  assign t[245] = t[300] ^ x[39];
  assign t[246] = t[301] ^ x[40];
  assign t[247] = t[302] ^ x[45];
  assign t[248] = t[303] ^ x[46];
  assign t[249] = t[304] ^ x[51];
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = t[305] ^ x[52];
  assign t[251] = t[306] ^ x[59];
  assign t[252] = t[307] ^ x[60];
  assign t[253] = t[308] ^ x[63];
  assign t[254] = t[309] ^ x[64];
  assign t[255] = t[310] ^ x[69];
  assign t[256] = t[311] ^ x[70];
  assign t[257] = t[312] ^ x[77];
  assign t[258] = t[313] ^ x[78];
  assign t[259] = t[314] ^ x[81];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[315] ^ x[82];
  assign t[261] = t[316] ^ x[83];
  assign t[262] = t[317] ^ x[84];
  assign t[263] = t[318] ^ x[85];
  assign t[264] = t[319] ^ x[86];
  assign t[265] = t[320] ^ x[87];
  assign t[266] = t[321] ^ x[88];
  assign t[267] = t[322] ^ x[89];
  assign t[268] = t[323] ^ x[90];
  assign t[269] = t[324] ^ x[95];
  assign t[26] = ~(t[41] & t[42]);
  assign t[270] = t[325] ^ x[96];
  assign t[271] = t[326] ^ x[97];
  assign t[272] = t[327] ^ x[98];
  assign t[273] = t[328] ^ x[103];
  assign t[274] = t[329] ^ x[104];
  assign t[275] = t[330] ^ x[105];
  assign t[276] = t[331] ^ x[106];
  assign t[277] = t[332] ^ x[107];
  assign t[278] = t[333] ^ x[108];
  assign t[279] = t[334] ^ x[109];
  assign t[27] = ~(t[43] & t[113]);
  assign t[280] = t[335] ^ x[110];
  assign t[281] = t[336] ^ x[111];
  assign t[282] = t[337] ^ x[112];
  assign t[283] = t[338] ^ x[113];
  assign t[284] = t[339] ^ x[114];
  assign t[285] = t[340] ^ x[115];
  assign t[286] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[287] = (x[2]);
  assign t[288] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[289] = (x[9]);
  assign t[28] = t[44] ? x[30] : x[29];
  assign t[290] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[291] = (x[12]);
  assign t[292] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[293] = (x[15]);
  assign t[294] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[295] = (x[18]);
  assign t[296] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[297] = (x[24]);
  assign t[298] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[299] = (x[32]);
  assign t[29] = ~(t[45] & t[46]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = (x[26]);
  assign t[301] = (x[23]);
  assign t[302] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[303] = (x[42]);
  assign t[304] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[305] = (x[48]);
  assign t[306] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[307] = (x[56]);
  assign t[308] = (x[34]);
  assign t[309] = (x[31]);
  assign t[30] = ~(t[47] & t[48]);
  assign t[310] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[311] = (x[66]);
  assign t[312] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[313] = (x[74]);
  assign t[314] = (x[25]);
  assign t[315] = (x[44]);
  assign t[316] = (x[41]);
  assign t[317] = (x[50]);
  assign t[318] = (x[47]);
  assign t[319] = (x[58]);
  assign t[31] = t[49] ^ t[37];
  assign t[320] = (x[55]);
  assign t[321] = (x[33]);
  assign t[322] = (x[68]);
  assign t[323] = (x[65]);
  assign t[324] = (x[91] & ~x[92] & ~x[93] & ~x[94]) | (~x[91] & x[92] & ~x[93] & ~x[94]) | (~x[91] & ~x[92] & x[93] & ~x[94]) | (~x[91] & ~x[92] & ~x[93] & x[94]) | (x[91] & x[92] & x[93] & ~x[94]) | (x[91] & x[92] & ~x[93] & x[94]) | (x[91] & ~x[92] & x[93] & x[94]) | (~x[91] & x[92] & x[93] & x[94]);
  assign t[325] = (x[92]);
  assign t[326] = (x[76]);
  assign t[327] = (x[73]);
  assign t[328] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[329] = (x[100]);
  assign t[32] = ~(t[50] & t[51]);
  assign t[330] = (x[43]);
  assign t[331] = (x[49]);
  assign t[332] = (x[57]);
  assign t[333] = (x[67]);
  assign t[334] = (x[94]);
  assign t[335] = (x[91]);
  assign t[336] = (x[75]);
  assign t[337] = (x[102]);
  assign t[338] = (x[99]);
  assign t[339] = (x[93]);
  assign t[33] = t[52] ^ t[30];
  assign t[340] = (x[101]);
  assign t[34] = ~(t[53] & t[54]);
  assign t[35] = ~(t[55] & t[114]);
  assign t[36] = t[111] ? x[38] : x[37];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = t[58] ^ t[59];
  assign t[39] = ~(t[60] & t[61]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[62] ^ t[63];
  assign t[41] = ~(t[115]);
  assign t[42] = ~(t[116]);
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = ~(t[66]);
  assign t[45] = ~(t[67] & t[68]);
  assign t[46] = ~(t[69] & t[117]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[118]);
  assign t[49] = t[44] ? x[54] : x[53];
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[119]);
  assign t[52] = t[111] ? x[62] : x[61];
  assign t[53] = ~(t[120]);
  assign t[54] = ~(t[121]);
  assign t[55] = ~(t[76] & t[77]);
  assign t[56] = ~(t[78] & t[79]);
  assign t[57] = ~(t[80] & t[122]);
  assign t[58] = t[111] ? x[72] : x[71];
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[123]);
  assign t[62] = t[44] ? x[80] : x[79];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[116] & t[115]);
  assign t[65] = ~(t[124]);
  assign t[66] = ~(t[111]);
  assign t[67] = ~(t[125]);
  assign t[68] = ~(t[126]);
  assign t[69] = ~(t[88] & t[89]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[128]);
  assign t[72] = ~(t[90] & t[91]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[92] & t[93]);
  assign t[76] = ~(t[121] & t[120]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = ~(t[109] & t[110]);
  assign t[80] = ~(t[94] & t[95]);
  assign t[81] = ~(t[96] & t[97]);
  assign t[82] = ~(t[98] & t[134]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[99] & t[100]);
  assign t[86] = ~(t[101] & t[102]);
  assign t[87] = ~(t[103] & t[137]);
  assign t[88] = ~(t[126] & t[125]);
  assign t[89] = ~(t[138]);
  assign t[8] = ~(t[111] & t[112]);
  assign t[90] = ~(t[128] & t[127]);
  assign t[91] = ~(t[139]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[140]);
  assign t[94] = ~(t[133] & t[132]);
  assign t[95] = ~(t[141]);
  assign t[96] = ~(t[142]);
  assign t[97] = ~(t[143]);
  assign t[98] = ~(t[104] & t[105]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [106:0] x;
 output y;

 wire [279:0] t;
  assign t[0] = t[1] ? t[2] : t[92];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = t[156] ^ x[5];
  assign t[125] = t[157] ^ x[11];
  assign t[126] = t[158] ^ x[14];
  assign t[127] = t[159] ^ x[17];
  assign t[128] = t[160] ^ x[20];
  assign t[129] = t[161] ^ x[28];
  assign t[12] = t[95] ? x[21] : x[22];
  assign t[130] = t[162] ^ x[29];
  assign t[131] = t[163] ^ x[37];
  assign t[132] = t[164] ^ x[38];
  assign t[133] = t[165] ^ x[41];
  assign t[134] = t[166] ^ x[47];
  assign t[135] = t[167] ^ x[48];
  assign t[136] = t[168] ^ x[54];
  assign t[137] = t[169] ^ x[55];
  assign t[138] = t[170] ^ x[63];
  assign t[139] = t[171] ^ x[64];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = t[172] ^ x[67];
  assign t[141] = t[173] ^ x[73];
  assign t[142] = t[174] ^ x[74];
  assign t[143] = t[175] ^ x[82];
  assign t[144] = t[176] ^ x[83];
  assign t[145] = t[177] ^ x[86];
  assign t[146] = t[178] ^ x[87];
  assign t[147] = t[179] ^ x[88];
  assign t[148] = t[180] ^ x[89];
  assign t[149] = t[181] ^ x[95];
  assign t[14] = x[7] ? t[19] : t[18];
  assign t[150] = t[182] ^ x[96];
  assign t[151] = t[183] ^ x[97];
  assign t[152] = t[184] ^ x[103];
  assign t[153] = t[185] ^ x[104];
  assign t[154] = t[186] ^ x[105];
  assign t[155] = t[187] ^ x[106];
  assign t[156] = (~t[188] & t[189]);
  assign t[157] = (~t[190] & t[191]);
  assign t[158] = (~t[192] & t[193]);
  assign t[159] = (~t[194] & t[195]);
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = (~t[196] & t[197]);
  assign t[161] = (~t[198] & t[199]);
  assign t[162] = (~t[198] & t[200]);
  assign t[163] = (~t[201] & t[202]);
  assign t[164] = (~t[201] & t[203]);
  assign t[165] = (~t[198] & t[204]);
  assign t[166] = (~t[205] & t[206]);
  assign t[167] = (~t[205] & t[207]);
  assign t[168] = (~t[208] & t[209]);
  assign t[169] = (~t[208] & t[210]);
  assign t[16] = x[7] ? t[23] : t[22];
  assign t[170] = (~t[211] & t[212]);
  assign t[171] = (~t[211] & t[213]);
  assign t[172] = (~t[201] & t[214]);
  assign t[173] = (~t[215] & t[216]);
  assign t[174] = (~t[215] & t[217]);
  assign t[175] = (~t[218] & t[219]);
  assign t[176] = (~t[218] & t[220]);
  assign t[177] = (~t[205] & t[221]);
  assign t[178] = (~t[208] & t[222]);
  assign t[179] = (~t[211] & t[223]);
  assign t[17] = ~(t[24] ^ t[25]);
  assign t[180] = (~t[215] & t[224]);
  assign t[181] = (~t[225] & t[226]);
  assign t[182] = (~t[225] & t[227]);
  assign t[183] = (~t[218] & t[228]);
  assign t[184] = (~t[229] & t[230]);
  assign t[185] = (~t[229] & t[231]);
  assign t[186] = (~t[225] & t[232]);
  assign t[187] = (~t[229] & t[233]);
  assign t[188] = t[234] ^ x[4];
  assign t[189] = t[235] ^ x[5];
  assign t[18] = ~(t[26] & t[27]);
  assign t[190] = t[236] ^ x[10];
  assign t[191] = t[237] ^ x[11];
  assign t[192] = t[238] ^ x[13];
  assign t[193] = t[239] ^ x[14];
  assign t[194] = t[240] ^ x[16];
  assign t[195] = t[241] ^ x[17];
  assign t[196] = t[242] ^ x[19];
  assign t[197] = t[243] ^ x[20];
  assign t[198] = t[244] ^ x[27];
  assign t[199] = t[245] ^ x[28];
  assign t[19] = t[28] ^ t[29];
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[246] ^ x[29];
  assign t[201] = t[247] ^ x[36];
  assign t[202] = t[248] ^ x[37];
  assign t[203] = t[249] ^ x[38];
  assign t[204] = t[250] ^ x[41];
  assign t[205] = t[251] ^ x[46];
  assign t[206] = t[252] ^ x[47];
  assign t[207] = t[253] ^ x[48];
  assign t[208] = t[254] ^ x[53];
  assign t[209] = t[255] ^ x[54];
  assign t[20] = x[7] ? t[31] : t[30];
  assign t[210] = t[256] ^ x[55];
  assign t[211] = t[257] ^ x[62];
  assign t[212] = t[258] ^ x[63];
  assign t[213] = t[259] ^ x[64];
  assign t[214] = t[260] ^ x[67];
  assign t[215] = t[261] ^ x[72];
  assign t[216] = t[262] ^ x[73];
  assign t[217] = t[263] ^ x[74];
  assign t[218] = t[264] ^ x[81];
  assign t[219] = t[265] ^ x[82];
  assign t[21] = x[7] ? t[33] : t[32];
  assign t[220] = t[266] ^ x[83];
  assign t[221] = t[267] ^ x[86];
  assign t[222] = t[268] ^ x[87];
  assign t[223] = t[269] ^ x[88];
  assign t[224] = t[270] ^ x[89];
  assign t[225] = t[271] ^ x[94];
  assign t[226] = t[272] ^ x[95];
  assign t[227] = t[273] ^ x[96];
  assign t[228] = t[274] ^ x[97];
  assign t[229] = t[275] ^ x[102];
  assign t[22] = ~(t[34] & t[35]);
  assign t[230] = t[276] ^ x[103];
  assign t[231] = t[277] ^ x[104];
  assign t[232] = t[278] ^ x[105];
  assign t[233] = t[279] ^ x[106];
  assign t[234] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[235] = (x[1]);
  assign t[236] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[237] = (x[9]);
  assign t[238] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[239] = (x[12]);
  assign t[23] = t[36] ^ t[22];
  assign t[240] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[241] = (x[15]);
  assign t[242] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[243] = (x[18]);
  assign t[244] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[245] = (x[25]);
  assign t[246] = (x[23]);
  assign t[247] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[248] = (x[34]);
  assign t[249] = (x[32]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = (x[26]);
  assign t[251] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[252] = (x[44]);
  assign t[253] = (x[42]);
  assign t[254] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[255] = (x[51]);
  assign t[256] = (x[49]);
  assign t[257] = (x[58] & ~x[59] & ~x[60] & ~x[61]) | (~x[58] & x[59] & ~x[60] & ~x[61]) | (~x[58] & ~x[59] & x[60] & ~x[61]) | (~x[58] & ~x[59] & ~x[60] & x[61]) | (x[58] & x[59] & x[60] & ~x[61]) | (x[58] & x[59] & ~x[60] & x[61]) | (x[58] & ~x[59] & x[60] & x[61]) | (~x[58] & x[59] & x[60] & x[61]);
  assign t[258] = (x[60]);
  assign t[259] = (x[58]);
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = (x[35]);
  assign t[261] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[262] = (x[70]);
  assign t[263] = (x[68]);
  assign t[264] = (x[77] & ~x[78] & ~x[79] & ~x[80]) | (~x[77] & x[78] & ~x[79] & ~x[80]) | (~x[77] & ~x[78] & x[79] & ~x[80]) | (~x[77] & ~x[78] & ~x[79] & x[80]) | (x[77] & x[78] & x[79] & ~x[80]) | (x[77] & x[78] & ~x[79] & x[80]) | (x[77] & ~x[78] & x[79] & x[80]) | (~x[77] & x[78] & x[79] & x[80]);
  assign t[265] = (x[79]);
  assign t[266] = (x[77]);
  assign t[267] = (x[45]);
  assign t[268] = (x[52]);
  assign t[269] = (x[61]);
  assign t[26] = ~(t[97] & t[41]);
  assign t[270] = (x[71]);
  assign t[271] = (x[90] & ~x[91] & ~x[92] & ~x[93]) | (~x[90] & x[91] & ~x[92] & ~x[93]) | (~x[90] & ~x[91] & x[92] & ~x[93]) | (~x[90] & ~x[91] & ~x[92] & x[93]) | (x[90] & x[91] & x[92] & ~x[93]) | (x[90] & x[91] & ~x[92] & x[93]) | (x[90] & ~x[91] & x[92] & x[93]) | (~x[90] & x[91] & x[92] & x[93]);
  assign t[272] = (x[92]);
  assign t[273] = (x[90]);
  assign t[274] = (x[80]);
  assign t[275] = (x[98] & ~x[99] & ~x[100] & ~x[101]) | (~x[98] & x[99] & ~x[100] & ~x[101]) | (~x[98] & ~x[99] & x[100] & ~x[101]) | (~x[98] & ~x[99] & ~x[100] & x[101]) | (x[98] & x[99] & x[100] & ~x[101]) | (x[98] & x[99] & ~x[100] & x[101]) | (x[98] & ~x[99] & x[100] & x[101]) | (~x[98] & x[99] & x[100] & x[101]);
  assign t[276] = (x[100]);
  assign t[277] = (x[98]);
  assign t[278] = (x[93]);
  assign t[279] = (x[101]);
  assign t[27] = ~(t[98] & t[42]);
  assign t[28] = t[43] ? x[31] : x[30];
  assign t[29] = ~(t[44] & t[45]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = ~(t[46] & t[47]);
  assign t[31] = t[48] ^ t[32];
  assign t[32] = ~(t[49] & t[50]);
  assign t[33] = t[51] ^ t[37];
  assign t[34] = ~(t[99] & t[52]);
  assign t[35] = ~(t[100] & t[53]);
  assign t[36] = t[95] ? x[40] : x[39];
  assign t[37] = ~(t[54] & t[55]);
  assign t[38] = t[56] ^ t[57];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[60] ^ t[61];
  assign t[41] = ~(t[101]);
  assign t[42] = ~(t[101] & t[62]);
  assign t[43] = ~(t[63]);
  assign t[44] = ~(t[102] & t[64]);
  assign t[45] = ~(t[103] & t[65]);
  assign t[46] = ~(t[104] & t[66]);
  assign t[47] = ~(t[105] & t[67]);
  assign t[48] = t[68] ? x[57] : x[56];
  assign t[49] = ~(t[106] & t[69]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[107] & t[70]);
  assign t[51] = t[71] ? x[66] : x[65];
  assign t[52] = ~(t[108]);
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = ~(t[109] & t[73]);
  assign t[55] = ~(t[110] & t[74]);
  assign t[56] = t[95] ? x[76] : x[75];
  assign t[57] = ~(t[75] & t[76]);
  assign t[58] = ~(t[111] & t[77]);
  assign t[59] = ~(t[112] & t[78]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[43] ? x[85] : x[84];
  assign t[61] = ~(t[79] & t[80]);
  assign t[62] = ~(t[97]);
  assign t[63] = ~(t[95]);
  assign t[64] = ~(t[113]);
  assign t[65] = ~(t[113] & t[81]);
  assign t[66] = ~(t[114]);
  assign t[67] = ~(t[114] & t[82]);
  assign t[68] = ~(t[63]);
  assign t[69] = ~(t[115]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[63]);
  assign t[72] = ~(t[99]);
  assign t[73] = ~(t[116]);
  assign t[74] = ~(t[116] & t[84]);
  assign t[75] = ~(t[117] & t[85]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119]);
  assign t[78] = ~(t[119] & t[87]);
  assign t[79] = ~(t[120] & t[88]);
  assign t[7] = ~(t[93] & t[94]);
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[102]);
  assign t[82] = ~(t[104]);
  assign t[83] = ~(t[106]);
  assign t[84] = ~(t[109]);
  assign t[85] = ~(t[122]);
  assign t[86] = ~(t[122] & t[90]);
  assign t[87] = ~(t[111]);
  assign t[88] = ~(t[123]);
  assign t[89] = ~(t[123] & t[91]);
  assign t[8] = ~(t[95] & t[96]);
  assign t[90] = ~(t[117]);
  assign t[91] = ~(t[120]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [115:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[224]);
  assign t[101] = ~(t[213] | t[214]);
  assign t[102] = ~(t[138] & t[140]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[226]);
  assign t[105] = ~(t[141] | t[142]);
  assign t[106] = ~(t[143] | t[144]);
  assign t[107] = ~(t[227] | t[145]);
  assign t[108] = t[204] ? x[94] : x[93];
  assign t[109] = ~(t[146] & t[147]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[228]);
  assign t[111] = ~(t[229]);
  assign t[112] = ~(t[148] | t[149]);
  assign t[113] = ~(t[150] | t[151]);
  assign t[114] = ~(t[230] | t[152]);
  assign t[115] = t[204] ? x[104] : x[103];
  assign t[116] = ~(t[146] & t[153]);
  assign t[117] = ~(t[122] | t[202]);
  assign t[118] = ~(t[154] & t[155]);
  assign t[119] = ~(t[203] | t[156]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = t[80] & t[202];
  assign t[121] = ~(t[122] | t[157]);
  assign t[122] = ~(t[204]);
  assign t[123] = t[202] ? t[159] : t[158];
  assign t[124] = ~(t[160] & t[205]);
  assign t[125] = ~(t[161] & t[156]);
  assign t[126] = ~(t[231]);
  assign t[127] = ~(t[218] | t[219]);
  assign t[128] = ~(t[162] & t[163]);
  assign t[129] = ~(t[164] & t[79]);
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = ~(t[80] | t[165]);
  assign t[131] = ~(t[80] | t[166]);
  assign t[132] = ~(t[232]);
  assign t[133] = ~(t[220] | t[221]);
  assign t[134] = ~(t[130] | t[167]);
  assign t[135] = ~(t[168] | t[169]);
  assign t[136] = ~(t[233]);
  assign t[137] = ~(t[222] | t[223]);
  assign t[138] = ~(t[49] | t[170]);
  assign t[139] = ~(t[171] | t[172]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = ~(t[167] | t[131]);
  assign t[141] = ~(t[234]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[235]);
  assign t[144] = ~(t[236]);
  assign t[145] = ~(t[173] | t[174]);
  assign t[146] = ~(t[49] | t[175]);
  assign t[147] = ~(t[121] | t[176]);
  assign t[148] = ~(t[237]);
  assign t[149] = ~(t[228] | t[229]);
  assign t[14] = x[7] ? t[21] : t[20];
  assign t[150] = ~(t[238]);
  assign t[151] = ~(t[239]);
  assign t[152] = ~(t[177] | t[178]);
  assign t[153] = ~(t[179] | t[131]);
  assign t[154] = ~(t[205] & t[180]);
  assign t[155] = ~(x[7] & t[119]);
  assign t[156] = ~(t[205]);
  assign t[157] = t[202] ? t[158] : t[159];
  assign t[158] = ~(t[180] & t[156]);
  assign t[159] = ~(x[7] & t[181]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = x[7] & t[203];
  assign t[161] = ~(x[7] | t[203]);
  assign t[162] = ~(t[171] | t[182]);
  assign t[163] = ~(t[122] & t[183]);
  assign t[164] = ~(t[184] & t[185]);
  assign t[165] = t[202] ? t[124] : t[125];
  assign t[166] = t[202] ? t[187] : t[186];
  assign t[167] = ~(t[80] | t[188]);
  assign t[168] = t[172] | t[189];
  assign t[169] = ~(t[190] & t[79]);
  assign t[16] = x[7] ? t[25] : t[24];
  assign t[170] = ~(t[80] | t[191]);
  assign t[171] = ~(t[122] | t[192]);
  assign t[172] = ~(t[193] & t[77]);
  assign t[173] = ~(t[240]);
  assign t[174] = ~(t[235] | t[236]);
  assign t[175] = ~(t[134] & t[164]);
  assign t[176] = t[170] | t[194];
  assign t[177] = ~(t[241]);
  assign t[178] = ~(t[238] | t[239]);
  assign t[179] = ~(t[80] | t[195]);
  assign t[17] = ~(t[26] ^ t[27]);
  assign t[180] = ~(x[7] | t[196]);
  assign t[181] = ~(t[203] | t[205]);
  assign t[182] = ~(t[80] | t[197]);
  assign t[183] = ~(t[159] & t[154]);
  assign t[184] = t[205] & t[117];
  assign t[185] = t[161] | t[160];
  assign t[186] = ~(t[161] & t[205]);
  assign t[187] = ~(t[160] & t[156]);
  assign t[188] = t[202] ? t[159] : t[154];
  assign t[189] = ~(t[80] | t[198]);
  assign t[18] = t[28] ? x[21] : x[22];
  assign t[190] = ~(t[194] | t[179]);
  assign t[191] = t[202] ? t[186] : t[187];
  assign t[192] = t[202] ? t[125] : t[187];
  assign t[193] = ~(t[199] | t[121]);
  assign t[194] = ~(t[76]);
  assign t[195] = t[202] ? t[155] : t[158];
  assign t[196] = ~(t[203]);
  assign t[197] = t[202] ? t[158] : t[155];
  assign t[198] = t[202] ? t[154] : t[159];
  assign t[199] = ~(t[122] | t[200]);
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[202] ? t[187] : t[125];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = ~(t[31] | t[32]);
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[33] ^ t[34]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = x[7] ? t[36] : t[35];
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = x[7] ? t[38] : t[37];
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[5];
  assign t[243] = t[284] ^ x[11];
  assign t[244] = t[285] ^ x[14];
  assign t[245] = t[286] ^ x[17];
  assign t[246] = t[287] ^ x[20];
  assign t[247] = t[288] ^ x[28];
  assign t[248] = t[289] ^ x[34];
  assign t[249] = t[290] ^ x[35];
  assign t[24] = ~(t[39] | t[40]);
  assign t[250] = t[291] ^ x[36];
  assign t[251] = t[292] ^ x[42];
  assign t[252] = t[293] ^ x[50];
  assign t[253] = t[294] ^ x[56];
  assign t[254] = t[295] ^ x[57];
  assign t[255] = t[296] ^ x[58];
  assign t[256] = t[297] ^ x[66];
  assign t[257] = t[298] ^ x[72];
  assign t[258] = t[299] ^ x[73];
  assign t[259] = t[300] ^ x[74];
  assign t[25] = ~(t[24] ^ t[41]);
  assign t[260] = t[301] ^ x[75];
  assign t[261] = t[302] ^ x[76];
  assign t[262] = t[303] ^ x[77];
  assign t[263] = t[304] ^ x[80];
  assign t[264] = t[305] ^ x[81];
  assign t[265] = t[306] ^ x[84];
  assign t[266] = t[307] ^ x[85];
  assign t[267] = t[308] ^ x[86];
  assign t[268] = t[309] ^ x[92];
  assign t[269] = t[310] ^ x[95];
  assign t[26] = x[7] ? t[43] : t[42];
  assign t[270] = t[311] ^ x[96];
  assign t[271] = t[312] ^ x[102];
  assign t[272] = t[313] ^ x[105];
  assign t[273] = t[314] ^ x[106];
  assign t[274] = t[315] ^ x[107];
  assign t[275] = t[316] ^ x[108];
  assign t[276] = t[317] ^ x[109];
  assign t[277] = t[318] ^ x[110];
  assign t[278] = t[319] ^ x[111];
  assign t[279] = t[320] ^ x[112];
  assign t[27] = x[7] ? t[45] : t[44];
  assign t[280] = t[321] ^ x[113];
  assign t[281] = t[322] ^ x[114];
  assign t[282] = t[323] ^ x[115];
  assign t[283] = (~t[324] & t[325]);
  assign t[284] = (~t[326] & t[327]);
  assign t[285] = (~t[328] & t[329]);
  assign t[286] = (~t[330] & t[331]);
  assign t[287] = (~t[332] & t[333]);
  assign t[288] = (~t[334] & t[335]);
  assign t[289] = (~t[336] & t[337]);
  assign t[28] = ~(t[46]);
  assign t[290] = (~t[334] & t[338]);
  assign t[291] = (~t[334] & t[339]);
  assign t[292] = (~t[340] & t[341]);
  assign t[293] = (~t[342] & t[343]);
  assign t[294] = (~t[344] & t[345]);
  assign t[295] = (~t[336] & t[346]);
  assign t[296] = (~t[336] & t[347]);
  assign t[297] = (~t[348] & t[349]);
  assign t[298] = (~t[350] & t[351]);
  assign t[299] = (~t[334] & t[352]);
  assign t[29] = ~(t[47] | t[48]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = (~t[340] & t[353]);
  assign t[301] = (~t[340] & t[354]);
  assign t[302] = (~t[342] & t[355]);
  assign t[303] = (~t[342] & t[356]);
  assign t[304] = (~t[344] & t[357]);
  assign t[305] = (~t[344] & t[358]);
  assign t[306] = (~t[336] & t[359]);
  assign t[307] = (~t[348] & t[360]);
  assign t[308] = (~t[348] & t[361]);
  assign t[309] = (~t[362] & t[363]);
  assign t[30] = ~(t[49]);
  assign t[310] = (~t[350] & t[364]);
  assign t[311] = (~t[350] & t[365]);
  assign t[312] = (~t[366] & t[367]);
  assign t[313] = (~t[340] & t[368]);
  assign t[314] = (~t[342] & t[369]);
  assign t[315] = (~t[344] & t[370]);
  assign t[316] = (~t[348] & t[371]);
  assign t[317] = (~t[362] & t[372]);
  assign t[318] = (~t[362] & t[373]);
  assign t[319] = (~t[350] & t[374]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (~t[366] & t[375]);
  assign t[321] = (~t[366] & t[376]);
  assign t[322] = (~t[362] & t[377]);
  assign t[323] = (~t[366] & t[378]);
  assign t[324] = t[379] ^ x[4];
  assign t[325] = t[380] ^ x[5];
  assign t[326] = t[381] ^ x[10];
  assign t[327] = t[382] ^ x[11];
  assign t[328] = t[383] ^ x[13];
  assign t[329] = t[384] ^ x[14];
  assign t[32] = ~(t[206] | t[52]);
  assign t[330] = t[385] ^ x[16];
  assign t[331] = t[386] ^ x[17];
  assign t[332] = t[387] ^ x[19];
  assign t[333] = t[388] ^ x[20];
  assign t[334] = t[389] ^ x[27];
  assign t[335] = t[390] ^ x[28];
  assign t[336] = t[391] ^ x[33];
  assign t[337] = t[392] ^ x[34];
  assign t[338] = t[393] ^ x[35];
  assign t[339] = t[394] ^ x[36];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[395] ^ x[41];
  assign t[341] = t[396] ^ x[42];
  assign t[342] = t[397] ^ x[49];
  assign t[343] = t[398] ^ x[50];
  assign t[344] = t[399] ^ x[55];
  assign t[345] = t[400] ^ x[56];
  assign t[346] = t[401] ^ x[57];
  assign t[347] = t[402] ^ x[58];
  assign t[348] = t[403] ^ x[65];
  assign t[349] = t[404] ^ x[66];
  assign t[34] = ~(t[55] ^ t[56]);
  assign t[350] = t[405] ^ x[71];
  assign t[351] = t[406] ^ x[72];
  assign t[352] = t[407] ^ x[73];
  assign t[353] = t[408] ^ x[74];
  assign t[354] = t[409] ^ x[75];
  assign t[355] = t[410] ^ x[76];
  assign t[356] = t[411] ^ x[77];
  assign t[357] = t[412] ^ x[80];
  assign t[358] = t[413] ^ x[81];
  assign t[359] = t[414] ^ x[84];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[415] ^ x[85];
  assign t[361] = t[416] ^ x[86];
  assign t[362] = t[417] ^ x[91];
  assign t[363] = t[418] ^ x[92];
  assign t[364] = t[419] ^ x[95];
  assign t[365] = t[420] ^ x[96];
  assign t[366] = t[421] ^ x[101];
  assign t[367] = t[422] ^ x[102];
  assign t[368] = t[423] ^ x[105];
  assign t[369] = t[424] ^ x[106];
  assign t[36] = ~(t[44] ^ t[59]);
  assign t[370] = t[425] ^ x[107];
  assign t[371] = t[426] ^ x[108];
  assign t[372] = t[427] ^ x[109];
  assign t[373] = t[428] ^ x[110];
  assign t[374] = t[429] ^ x[111];
  assign t[375] = t[430] ^ x[112];
  assign t[376] = t[431] ^ x[113];
  assign t[377] = t[432] ^ x[114];
  assign t[378] = t[433] ^ x[115];
  assign t[379] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = (x[0]);
  assign t[381] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[382] = (x[9]);
  assign t[383] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[384] = (x[12]);
  assign t[385] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[386] = (x[15]);
  assign t[387] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[388] = (x[18]);
  assign t[389] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[38] = ~(t[35] ^ t[62]);
  assign t[390] = (x[24]);
  assign t[391] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[392] = (x[30]);
  assign t[393] = (x[25]);
  assign t[394] = (x[26]);
  assign t[395] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[396] = (x[38]);
  assign t[397] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[398] = (x[46]);
  assign t[399] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[400] = (x[52]);
  assign t[401] = (x[31]);
  assign t[402] = (x[32]);
  assign t[403] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[404] = (x[62]);
  assign t[405] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[406] = (x[68]);
  assign t[407] = (x[23]);
  assign t[408] = (x[39]);
  assign t[409] = (x[40]);
  assign t[40] = ~(t[207] | t[65]);
  assign t[410] = (x[47]);
  assign t[411] = (x[48]);
  assign t[412] = (x[53]);
  assign t[413] = (x[54]);
  assign t[414] = (x[29]);
  assign t[415] = (x[63]);
  assign t[416] = (x[64]);
  assign t[417] = (x[87] & ~x[88] & ~x[89] & ~x[90]) | (~x[87] & x[88] & ~x[89] & ~x[90]) | (~x[87] & ~x[88] & x[89] & ~x[90]) | (~x[87] & ~x[88] & ~x[89] & x[90]) | (x[87] & x[88] & x[89] & ~x[90]) | (x[87] & x[88] & ~x[89] & x[90]) | (x[87] & ~x[88] & x[89] & x[90]) | (~x[87] & x[88] & x[89] & x[90]);
  assign t[418] = (x[88]);
  assign t[419] = (x[69]);
  assign t[41] = ~(t[66] ^ t[67]);
  assign t[420] = (x[70]);
  assign t[421] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[422] = (x[98]);
  assign t[423] = (x[37]);
  assign t[424] = (x[45]);
  assign t[425] = (x[51]);
  assign t[426] = (x[61]);
  assign t[427] = (x[89]);
  assign t[428] = (x[90]);
  assign t[429] = (x[67]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[99]);
  assign t[431] = (x[100]);
  assign t[432] = (x[87]);
  assign t[433] = (x[97]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[46] = ~(t[204]);
  assign t[47] = ~(t[76] & t[77]);
  assign t[48] = ~(t[78] & t[79]);
  assign t[49] = ~(t[80] | t[81]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[208]);
  assign t[51] = ~(t[209]);
  assign t[52] = ~(t[82] | t[83]);
  assign t[53] = ~(t[84] | t[85]);
  assign t[54] = ~(t[210] | t[86]);
  assign t[55] = t[87] ? x[44] : x[43];
  assign t[56] = ~(t[88] & t[89]);
  assign t[57] = ~(t[90] | t[91]);
  assign t[58] = ~(t[211] | t[92]);
  assign t[59] = ~(t[93] ^ t[94]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[95] | t[96]);
  assign t[61] = ~(t[212] | t[97]);
  assign t[62] = ~(t[98] ^ t[99]);
  assign t[63] = ~(t[213]);
  assign t[64] = ~(t[214]);
  assign t[65] = ~(t[100] | t[101]);
  assign t[66] = t[204] ? x[60] : x[59];
  assign t[67] = t[47] | t[102];
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = ~(t[215] | t[105]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[106] | t[107]);
  assign t[71] = ~(t[108] ^ t[109]);
  assign t[72] = ~(t[110] | t[111]);
  assign t[73] = ~(t[216] | t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[115] ^ t[116]);
  assign t[76] = ~(t[117] & t[118]);
  assign t[77] = ~(t[119] & t[120]);
  assign t[78] = ~(t[121]);
  assign t[79] = t[122] | t[123];
  assign t[7] = ~(t[202] & t[203]);
  assign t[80] = ~(t[122]);
  assign t[81] = t[202] ? t[125] : t[124];
  assign t[82] = ~(t[217]);
  assign t[83] = ~(t[208] | t[209]);
  assign t[84] = ~(t[218]);
  assign t[85] = ~(t[219]);
  assign t[86] = ~(t[126] | t[127]);
  assign t[87] = ~(t[46]);
  assign t[88] = ~(t[128] | t[129]);
  assign t[89] = ~(t[130] | t[131]);
  assign t[8] = ~(t[204] & t[205]);
  assign t[90] = ~(t[220]);
  assign t[91] = ~(t[221]);
  assign t[92] = ~(t[132] | t[133]);
  assign t[93] = t[87] ? x[79] : x[78];
  assign t[94] = ~(t[134] & t[135]);
  assign t[95] = ~(t[222]);
  assign t[96] = ~(t[223]);
  assign t[97] = ~(t[136] | t[137]);
  assign t[98] = t[87] ? x[83] : x[82];
  assign t[99] = ~(t[138] & t[139]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [172:0] x;
 output y;

 wire [672:0] t;
  assign t[0] = t[1] ? t[2] : t[403];
  assign t[100] = t[144] | t[145];
  assign t[101] = ~(t[425]);
  assign t[102] = ~(t[426]);
  assign t[103] = ~(t[146] | t[147]);
  assign t[104] = ~(t[148] | t[149]);
  assign t[105] = ~(t[427] | t[150]);
  assign t[106] = t[143] ? x[95] : x[94];
  assign t[107] = ~(t[151] & t[152]);
  assign t[108] = ~(t[428]);
  assign t[109] = ~(t[415] | t[416]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[429]);
  assign t[111] = ~(t[430]);
  assign t[112] = ~(t[153] | t[154]);
  assign t[113] = ~(t[155] | t[156]);
  assign t[114] = ~(t[431]);
  assign t[115] = ~(t[432]);
  assign t[116] = ~(t[157] | t[158]);
  assign t[117] = ~(t[159] | t[160]);
  assign t[118] = ~(t[433] | t[161]);
  assign t[119] = t[30] ? x[108] : x[107];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[162] & t[163]);
  assign t[121] = ~(t[434]);
  assign t[122] = ~(t[435]);
  assign t[123] = ~(t[164] | t[165]);
  assign t[124] = t[30] ? x[112] : x[111];
  assign t[125] = ~(t[166] & t[167]);
  assign t[126] = ~(t[128] | t[168]);
  assign t[127] = ~(t[86] | t[169]);
  assign t[128] = ~(t[406]);
  assign t[129] = ~(t[170] & t[171]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[407] & t[172];
  assign t[131] = t[173] | t[174];
  assign t[132] = t[404] ? t[170] : t[175];
  assign t[133] = ~(t[173] & t[176]);
  assign t[134] = ~(t[174] & t[407]);
  assign t[135] = ~(t[173] & t[407]);
  assign t[136] = ~(t[174] & t[176]);
  assign t[137] = ~(t[436]);
  assign t[138] = ~(t[421] | t[422]);
  assign t[139] = ~(t[405] | t[176]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[86] & t[404];
  assign t[141] = ~(t[437]);
  assign t[142] = ~(t[423] | t[424]);
  assign t[143] = ~(t[49]);
  assign t[144] = ~(t[177] & t[95]);
  assign t[145] = ~(t[86] | t[178]);
  assign t[146] = ~(t[438]);
  assign t[147] = ~(t[425] | t[426]);
  assign t[148] = ~(t[439]);
  assign t[149] = ~(t[440]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[179] | t[180]);
  assign t[151] = ~(t[52]);
  assign t[152] = ~(t[181] | t[145]);
  assign t[153] = ~(t[441]);
  assign t[154] = ~(t[429] | t[430]);
  assign t[155] = ~(t[86] | t[182]);
  assign t[156] = ~(t[32] & t[85]);
  assign t[157] = ~(t[442]);
  assign t[158] = ~(t[431] | t[432]);
  assign t[159] = ~(t[443]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[444]);
  assign t[161] = ~(t[183] | t[184]);
  assign t[162] = ~(t[52] | t[185]);
  assign t[163] = ~(t[100] | t[186]);
  assign t[164] = ~(t[445]);
  assign t[165] = ~(t[434] | t[435]);
  assign t[166] = ~(t[187] | t[155]);
  assign t[167] = ~(t[126] | t[144]);
  assign t[168] = t[404] ? t[133] : t[136];
  assign t[169] = t[404] ? t[175] : t[188];
  assign t[16] = ~(t[404] & t[405]);
  assign t[170] = ~(x[7] & t[189]);
  assign t[171] = ~(t[407] & t[190]);
  assign t[172] = ~(t[128] | t[404]);
  assign t[173] = ~(x[7] | t[405]);
  assign t[174] = x[7] & t[405];
  assign t[175] = ~(t[190] & t[176]);
  assign t[176] = ~(t[407]);
  assign t[177] = ~(t[191] | t[192]);
  assign t[178] = t[404] ? t[171] : t[170];
  assign t[179] = ~(t[446]);
  assign t[17] = ~(t[406] & t[407]);
  assign t[180] = ~(t[439] | t[440]);
  assign t[181] = ~(t[193]);
  assign t[182] = t[404] ? t[135] : t[136];
  assign t[183] = ~(t[447]);
  assign t[184] = ~(t[443] | t[444]);
  assign t[185] = ~(t[86] | t[194]);
  assign t[186] = ~(t[195] & t[85]);
  assign t[187] = ~(t[86] | t[196]);
  assign t[188] = ~(x[7] & t[139]);
  assign t[189] = ~(t[405] | t[407]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(x[7] | t[197]);
  assign t[191] = ~(t[128] | t[198]);
  assign t[192] = ~(t[128] | t[199]);
  assign t[193] = ~(t[200] | t[53]);
  assign t[194] = t[404] ? t[170] : t[171];
  assign t[195] = ~(t[201] | t[200]);
  assign t[196] = t[404] ? t[133] : t[134];
  assign t[197] = ~(t[405]);
  assign t[198] = t[404] ? t[136] : t[133];
  assign t[199] = t[404] ? t[175] : t[170];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[86] | t[202]);
  assign t[201] = ~(t[203]);
  assign t[202] = t[404] ? t[188] : t[175];
  assign t[203] = ~(t[172] & t[204]);
  assign t[204] = ~(t[171] & t[188]);
  assign t[205] = t[1] ? t[206] : t[448];
  assign t[206] = x[6] ? t[208] : t[207];
  assign t[207] = x[7] ? t[210] : t[209];
  assign t[208] = t[211] ^ x[126];
  assign t[209] = t[212] ^ t[213];
  assign t[20] = t[30] ? x[9] : x[10];
  assign t[210] = ~(t[214] ^ t[215]);
  assign t[211] = x[127] ^ x[128];
  assign t[212] = t[216] ? x[127] : x[128];
  assign t[213] = ~(t[217] ^ t[218]);
  assign t[214] = x[7] ? t[220] : t[219];
  assign t[215] = ~(t[221] ^ t[222]);
  assign t[216] = ~(t[49]);
  assign t[217] = x[7] ? t[224] : t[223];
  assign t[218] = ~(t[225] ^ t[226]);
  assign t[219] = ~(t[227] & t[228]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = t[229] ^ t[230];
  assign t[221] = x[7] ? t[232] : t[231];
  assign t[222] = x[7] ? t[234] : t[233];
  assign t[223] = ~(t[235] & t[236]);
  assign t[224] = t[237] ^ t[238];
  assign t[225] = x[7] ? t[240] : t[239];
  assign t[226] = x[7] ? t[242] : t[241];
  assign t[227] = ~(t[410] & t[55]);
  assign t[228] = ~(t[420] & t[243]);
  assign t[229] = t[30] ? x[130] : x[129];
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = ~(t[244] & t[245]);
  assign t[231] = ~(t[246] & t[247]);
  assign t[232] = t[248] ^ t[249];
  assign t[233] = ~(t[250] & t[251]);
  assign t[234] = t[252] ^ t[231];
  assign t[235] = ~(t[415] & t[69]);
  assign t[236] = ~(t[428] & t[253]);
  assign t[237] = t[30] ? x[132] : x[131];
  assign t[238] = ~(t[254] & t[255]);
  assign t[239] = ~(t[256] & t[257]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = t[258] ^ t[241];
  assign t[241] = ~(t[259] & t[260]);
  assign t[242] = t[261] ^ t[262];
  assign t[243] = ~(t[411] & t[54]);
  assign t[244] = ~(t[421] & t[92]);
  assign t[245] = ~(t[436] & t[263]);
  assign t[246] = ~(t[425] & t[102]);
  assign t[247] = ~(t[438] & t[264]);
  assign t[248] = t[143] ? x[134] : x[133];
  assign t[249] = ~(t[265] & t[266]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = ~(t[423] & t[97]);
  assign t[251] = ~(t[437] & t[267]);
  assign t[252] = t[143] ? x[136] : x[135];
  assign t[253] = ~(t[416] & t[68]);
  assign t[254] = ~(t[429] & t[111]);
  assign t[255] = ~(t[441] & t[268]);
  assign t[256] = ~(t[434] & t[122]);
  assign t[257] = ~(t[445] & t[269]);
  assign t[258] = t[143] ? x[138] : x[137];
  assign t[259] = ~(t[431] & t[115]);
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = ~(t[442] & t[270]);
  assign t[261] = t[30] ? x[140] : x[139];
  assign t[262] = ~(t[271] & t[272]);
  assign t[263] = ~(t[422] & t[91]);
  assign t[264] = ~(t[426] & t[101]);
  assign t[265] = ~(t[439] & t[149]);
  assign t[266] = ~(t[446] & t[273]);
  assign t[267] = ~(t[424] & t[96]);
  assign t[268] = ~(t[430] & t[110]);
  assign t[269] = ~(t[435] & t[121]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = ~(t[432] & t[114]);
  assign t[271] = ~(t[443] & t[160]);
  assign t[272] = ~(t[447] & t[274]);
  assign t[273] = ~(t[440] & t[148]);
  assign t[274] = ~(t[444] & t[159]);
  assign t[275] = t[1] ? t[276] : t[449];
  assign t[276] = x[6] ? t[278] : t[277];
  assign t[277] = x[7] ? t[280] : t[279];
  assign t[278] = t[281] ^ x[142];
  assign t[279] = t[282] ^ t[283];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = ~(t[284] ^ t[285]);
  assign t[281] = x[143] ^ x[144];
  assign t[282] = t[30] ? x[143] : x[144];
  assign t[283] = ~(t[286] ^ t[287]);
  assign t[284] = x[7] ? t[289] : t[288];
  assign t[285] = ~(t[290] ^ t[291]);
  assign t[286] = x[7] ? t[293] : t[292];
  assign t[287] = ~(t[294] ^ t[295]);
  assign t[288] = ~(t[296] & t[297]);
  assign t[289] = t[298] ^ t[299];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = x[7] ? t[301] : t[300];
  assign t[291] = x[7] ? t[303] : t[302];
  assign t[292] = ~(t[304] & t[305]);
  assign t[293] = t[306] ^ t[307];
  assign t[294] = x[7] ? t[309] : t[308];
  assign t[295] = x[7] ? t[311] : t[310];
  assign t[296] = ~(t[55] & t[89]);
  assign t[297] = ~(t[312] & t[408]);
  assign t[298] = t[30] ? x[146] : x[145];
  assign t[299] = ~(t[313] & t[314]);
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = ~(t[315] & t[316]);
  assign t[301] = t[317] ^ t[302];
  assign t[302] = ~(t[318] & t[319]);
  assign t[303] = t[320] ^ t[321];
  assign t[304] = ~(t[69] & t[108]);
  assign t[305] = ~(t[322] & t[409]);
  assign t[306] = t[143] ? x[148] : x[147];
  assign t[307] = ~(t[323] & t[324]);
  assign t[308] = ~(t[325] & t[326]);
  assign t[309] = t[327] ^ t[328];
  assign t[30] = ~(t[49]);
  assign t[310] = ~(t[329] & t[330]);
  assign t[311] = t[331] ^ t[308];
  assign t[312] = ~(t[332] & t[54]);
  assign t[313] = ~(t[92] & t[137]);
  assign t[314] = ~(t[333] & t[412]);
  assign t[315] = ~(t[97] & t[141]);
  assign t[316] = ~(t[334] & t[413]);
  assign t[317] = t[143] ? x[150] : x[149];
  assign t[318] = ~(t[102] & t[146]);
  assign t[319] = ~(t[335] & t[414]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = t[143] ? x[152] : x[151];
  assign t[321] = ~(t[336] & t[337]);
  assign t[322] = ~(t[338] & t[68]);
  assign t[323] = ~(t[111] & t[153]);
  assign t[324] = ~(t[339] & t[417]);
  assign t[325] = ~(t[115] & t[157]);
  assign t[326] = ~(t[340] & t[418]);
  assign t[327] = t[30] ? x[154] : x[153];
  assign t[328] = ~(t[341] & t[342]);
  assign t[329] = ~(t[122] & t[164]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = ~(t[343] & t[419]);
  assign t[331] = t[406] ? x[156] : x[155];
  assign t[332] = ~(t[420] & t[411]);
  assign t[333] = ~(t[344] & t[91]);
  assign t[334] = ~(t[345] & t[96]);
  assign t[335] = ~(t[346] & t[101]);
  assign t[336] = ~(t[149] & t[179]);
  assign t[337] = ~(t[347] & t[427]);
  assign t[338] = ~(t[428] & t[416]);
  assign t[339] = ~(t[348] & t[110]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = ~(t[349] & t[114]);
  assign t[341] = ~(t[160] & t[183]);
  assign t[342] = ~(t[350] & t[433]);
  assign t[343] = ~(t[351] & t[121]);
  assign t[344] = ~(t[436] & t[422]);
  assign t[345] = ~(t[437] & t[424]);
  assign t[346] = ~(t[438] & t[426]);
  assign t[347] = ~(t[352] & t[148]);
  assign t[348] = ~(t[441] & t[430]);
  assign t[349] = ~(t[442] & t[432]);
  assign t[34] = ~(t[408] | t[56]);
  assign t[350] = ~(t[353] & t[159]);
  assign t[351] = ~(t[445] & t[435]);
  assign t[352] = ~(t[446] & t[440]);
  assign t[353] = ~(t[447] & t[444]);
  assign t[354] = t[1] ? t[355] : t[450];
  assign t[355] = x[6] ? t[357] : t[356];
  assign t[356] = x[7] ? t[359] : t[358];
  assign t[357] = t[360] ^ x[158];
  assign t[358] = t[361] ^ t[362];
  assign t[359] = ~(t[363] ^ t[364]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = x[159] ^ x[160];
  assign t[361] = t[30] ? x[159] : x[160];
  assign t[362] = ~(t[365] ^ t[366]);
  assign t[363] = x[7] ? t[368] : t[367];
  assign t[364] = ~(t[369] ^ t[370]);
  assign t[365] = x[7] ? t[372] : t[371];
  assign t[366] = ~(t[373] ^ t[374]);
  assign t[367] = ~(t[296] & t[375]);
  assign t[368] = t[376] ^ t[377];
  assign t[369] = x[7] ? t[379] : t[378];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = x[7] ? t[381] : t[380];
  assign t[371] = ~(t[304] & t[382]);
  assign t[372] = t[383] ^ t[384];
  assign t[373] = x[7] ? t[386] : t[385];
  assign t[374] = x[7] ? t[388] : t[387];
  assign t[375] = t[33] | t[408];
  assign t[376] = t[30] ? x[162] : x[161];
  assign t[377] = ~(t[313] & t[389]);
  assign t[378] = ~(t[315] & t[390]);
  assign t[379] = t[391] ^ t[380];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = ~(t[318] & t[392]);
  assign t[381] = t[393] ^ t[394];
  assign t[382] = t[41] | t[409];
  assign t[383] = t[216] ? x[164] : x[163];
  assign t[384] = ~(t[323] & t[395]);
  assign t[385] = ~(t[325] & t[396]);
  assign t[386] = t[397] ^ t[398];
  assign t[387] = ~(t[329] & t[399]);
  assign t[388] = t[400] ^ t[385];
  assign t[389] = t[57] | t[412];
  assign t[38] = ~(t[39] ^ t[63]);
  assign t[390] = t[61] | t[413];
  assign t[391] = t[143] ? x[166] : x[165];
  assign t[392] = t[64] | t[414];
  assign t[393] = t[143] ? x[168] : x[167];
  assign t[394] = ~(t[336] & t[401]);
  assign t[395] = t[71] | t[417];
  assign t[396] = t[75] | t[418];
  assign t[397] = t[30] ? x[170] : x[169];
  assign t[398] = ~(t[341] & t[402]);
  assign t[399] = t[79] | t[419];
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[30] ? x[172] : x[171];
  assign t[401] = t[104] | t[427];
  assign t[402] = t[117] | t[433];
  assign t[403] = (t[451]);
  assign t[404] = (t[452]);
  assign t[405] = (t[453]);
  assign t[406] = (t[454]);
  assign t[407] = (t[455]);
  assign t[408] = (t[456]);
  assign t[409] = (t[457]);
  assign t[40] = ~(t[66] ^ t[67]);
  assign t[410] = (t[458]);
  assign t[411] = (t[459]);
  assign t[412] = (t[460]);
  assign t[413] = (t[461]);
  assign t[414] = (t[462]);
  assign t[415] = (t[463]);
  assign t[416] = (t[464]);
  assign t[417] = (t[465]);
  assign t[418] = (t[466]);
  assign t[419] = (t[467]);
  assign t[41] = ~(t[68] | t[69]);
  assign t[420] = (t[468]);
  assign t[421] = (t[469]);
  assign t[422] = (t[470]);
  assign t[423] = (t[471]);
  assign t[424] = (t[472]);
  assign t[425] = (t[473]);
  assign t[426] = (t[474]);
  assign t[427] = (t[475]);
  assign t[428] = (t[476]);
  assign t[429] = (t[477]);
  assign t[42] = ~(t[409] | t[70]);
  assign t[430] = (t[478]);
  assign t[431] = (t[479]);
  assign t[432] = (t[480]);
  assign t[433] = (t[481]);
  assign t[434] = (t[482]);
  assign t[435] = (t[483]);
  assign t[436] = (t[484]);
  assign t[437] = (t[485]);
  assign t[438] = (t[486]);
  assign t[439] = (t[487]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[440] = (t[488]);
  assign t[441] = (t[489]);
  assign t[442] = (t[490]);
  assign t[443] = (t[491]);
  assign t[444] = (t[492]);
  assign t[445] = (t[493]);
  assign t[446] = (t[494]);
  assign t[447] = (t[495]);
  assign t[448] = (t[496]);
  assign t[449] = (t[497]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[450] = (t[498]);
  assign t[451] = t[499] ^ x[5];
  assign t[452] = t[500] ^ x[13];
  assign t[453] = t[501] ^ x[16];
  assign t[454] = t[502] ^ x[19];
  assign t[455] = t[503] ^ x[22];
  assign t[456] = t[504] ^ x[28];
  assign t[457] = t[505] ^ x[34];
  assign t[458] = t[506] ^ x[35];
  assign t[459] = t[507] ^ x[36];
  assign t[45] = ~(t[75] | t[76]);
  assign t[460] = t[508] ^ x[42];
  assign t[461] = t[509] ^ x[50];
  assign t[462] = t[510] ^ x[56];
  assign t[463] = t[511] ^ x[57];
  assign t[464] = t[512] ^ x[58];
  assign t[465] = t[513] ^ x[64];
  assign t[466] = t[514] ^ x[72];
  assign t[467] = t[515] ^ x[78];
  assign t[468] = t[516] ^ x[79];
  assign t[469] = t[517] ^ x[80];
  assign t[46] = ~(t[77] ^ t[78]);
  assign t[470] = t[518] ^ x[81];
  assign t[471] = t[519] ^ x[82];
  assign t[472] = t[520] ^ x[83];
  assign t[473] = t[521] ^ x[86];
  assign t[474] = t[522] ^ x[87];
  assign t[475] = t[523] ^ x[93];
  assign t[476] = t[524] ^ x[96];
  assign t[477] = t[525] ^ x[97];
  assign t[478] = t[526] ^ x[98];
  assign t[479] = t[527] ^ x[99];
  assign t[47] = ~(t[79] | t[80]);
  assign t[480] = t[528] ^ x[100];
  assign t[481] = t[529] ^ x[106];
  assign t[482] = t[530] ^ x[109];
  assign t[483] = t[531] ^ x[110];
  assign t[484] = t[532] ^ x[113];
  assign t[485] = t[533] ^ x[114];
  assign t[486] = t[534] ^ x[115];
  assign t[487] = t[535] ^ x[116];
  assign t[488] = t[536] ^ x[117];
  assign t[489] = t[537] ^ x[118];
  assign t[48] = ~(t[45] ^ t[81]);
  assign t[490] = t[538] ^ x[119];
  assign t[491] = t[539] ^ x[120];
  assign t[492] = t[540] ^ x[121];
  assign t[493] = t[541] ^ x[122];
  assign t[494] = t[542] ^ x[123];
  assign t[495] = t[543] ^ x[124];
  assign t[496] = t[544] ^ x[125];
  assign t[497] = t[545] ^ x[141];
  assign t[498] = t[546] ^ x[157];
  assign t[499] = (~t[547] & t[548]);
  assign t[49] = ~(t[406]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[549] & t[550]);
  assign t[501] = (~t[551] & t[552]);
  assign t[502] = (~t[553] & t[554]);
  assign t[503] = (~t[555] & t[556]);
  assign t[504] = (~t[557] & t[558]);
  assign t[505] = (~t[559] & t[560]);
  assign t[506] = (~t[557] & t[561]);
  assign t[507] = (~t[557] & t[562]);
  assign t[508] = (~t[563] & t[564]);
  assign t[509] = (~t[565] & t[566]);
  assign t[50] = ~(t[82] & t[83]);
  assign t[510] = (~t[567] & t[568]);
  assign t[511] = (~t[559] & t[569]);
  assign t[512] = (~t[559] & t[570]);
  assign t[513] = (~t[571] & t[572]);
  assign t[514] = (~t[573] & t[574]);
  assign t[515] = (~t[575] & t[576]);
  assign t[516] = (~t[557] & t[577]);
  assign t[517] = (~t[563] & t[578]);
  assign t[518] = (~t[563] & t[579]);
  assign t[519] = (~t[565] & t[580]);
  assign t[51] = ~(t[84] & t[85]);
  assign t[520] = (~t[565] & t[581]);
  assign t[521] = (~t[567] & t[582]);
  assign t[522] = (~t[567] & t[583]);
  assign t[523] = (~t[584] & t[585]);
  assign t[524] = (~t[559] & t[586]);
  assign t[525] = (~t[571] & t[587]);
  assign t[526] = (~t[571] & t[588]);
  assign t[527] = (~t[573] & t[589]);
  assign t[528] = (~t[573] & t[590]);
  assign t[529] = (~t[591] & t[592]);
  assign t[52] = ~(t[86] | t[87]);
  assign t[530] = (~t[575] & t[593]);
  assign t[531] = (~t[575] & t[594]);
  assign t[532] = (~t[563] & t[595]);
  assign t[533] = (~t[565] & t[596]);
  assign t[534] = (~t[567] & t[597]);
  assign t[535] = (~t[584] & t[598]);
  assign t[536] = (~t[584] & t[599]);
  assign t[537] = (~t[571] & t[600]);
  assign t[538] = (~t[573] & t[601]);
  assign t[539] = (~t[591] & t[602]);
  assign t[53] = ~(t[86] | t[88]);
  assign t[540] = (~t[591] & t[603]);
  assign t[541] = (~t[575] & t[604]);
  assign t[542] = (~t[584] & t[605]);
  assign t[543] = (~t[591] & t[606]);
  assign t[544] = (~t[547] & t[607]);
  assign t[545] = (~t[547] & t[608]);
  assign t[546] = (~t[547] & t[609]);
  assign t[547] = t[610] ^ x[4];
  assign t[548] = t[611] ^ x[5];
  assign t[549] = t[612] ^ x[12];
  assign t[54] = ~(t[410]);
  assign t[550] = t[613] ^ x[13];
  assign t[551] = t[614] ^ x[15];
  assign t[552] = t[615] ^ x[16];
  assign t[553] = t[616] ^ x[18];
  assign t[554] = t[617] ^ x[19];
  assign t[555] = t[618] ^ x[21];
  assign t[556] = t[619] ^ x[22];
  assign t[557] = t[620] ^ x[27];
  assign t[558] = t[621] ^ x[28];
  assign t[559] = t[622] ^ x[33];
  assign t[55] = ~(t[411]);
  assign t[560] = t[623] ^ x[34];
  assign t[561] = t[624] ^ x[35];
  assign t[562] = t[625] ^ x[36];
  assign t[563] = t[626] ^ x[41];
  assign t[564] = t[627] ^ x[42];
  assign t[565] = t[628] ^ x[49];
  assign t[566] = t[629] ^ x[50];
  assign t[567] = t[630] ^ x[55];
  assign t[568] = t[631] ^ x[56];
  assign t[569] = t[632] ^ x[57];
  assign t[56] = ~(t[89] | t[90]);
  assign t[570] = t[633] ^ x[58];
  assign t[571] = t[634] ^ x[63];
  assign t[572] = t[635] ^ x[64];
  assign t[573] = t[636] ^ x[71];
  assign t[574] = t[637] ^ x[72];
  assign t[575] = t[638] ^ x[77];
  assign t[576] = t[639] ^ x[78];
  assign t[577] = t[640] ^ x[79];
  assign t[578] = t[641] ^ x[80];
  assign t[579] = t[642] ^ x[81];
  assign t[57] = ~(t[91] | t[92]);
  assign t[580] = t[643] ^ x[82];
  assign t[581] = t[644] ^ x[83];
  assign t[582] = t[645] ^ x[86];
  assign t[583] = t[646] ^ x[87];
  assign t[584] = t[647] ^ x[92];
  assign t[585] = t[648] ^ x[93];
  assign t[586] = t[649] ^ x[96];
  assign t[587] = t[650] ^ x[97];
  assign t[588] = t[651] ^ x[98];
  assign t[589] = t[652] ^ x[99];
  assign t[58] = ~(t[412] | t[93]);
  assign t[590] = t[653] ^ x[100];
  assign t[591] = t[654] ^ x[105];
  assign t[592] = t[655] ^ x[106];
  assign t[593] = t[656] ^ x[109];
  assign t[594] = t[657] ^ x[110];
  assign t[595] = t[658] ^ x[113];
  assign t[596] = t[659] ^ x[114];
  assign t[597] = t[660] ^ x[115];
  assign t[598] = t[661] ^ x[116];
  assign t[599] = t[662] ^ x[117];
  assign t[59] = t[30] ? x[44] : x[43];
  assign t[5] = t[9] ^ x[8];
  assign t[600] = t[663] ^ x[118];
  assign t[601] = t[664] ^ x[119];
  assign t[602] = t[665] ^ x[120];
  assign t[603] = t[666] ^ x[121];
  assign t[604] = t[667] ^ x[122];
  assign t[605] = t[668] ^ x[123];
  assign t[606] = t[669] ^ x[124];
  assign t[607] = t[670] ^ x[125];
  assign t[608] = t[671] ^ x[141];
  assign t[609] = t[672] ^ x[157];
  assign t[60] = ~(t[94] & t[95]);
  assign t[610] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[611] = (x[0]);
  assign t[612] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[613] = (x[11]);
  assign t[614] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[615] = (x[14]);
  assign t[616] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[617] = (x[17]);
  assign t[618] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[619] = (x[20]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[620] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[621] = (x[24]);
  assign t[622] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[623] = (x[30]);
  assign t[624] = (x[25]);
  assign t[625] = (x[26]);
  assign t[626] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[627] = (x[38]);
  assign t[628] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[629] = (x[46]);
  assign t[62] = ~(t[413] | t[98]);
  assign t[630] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[631] = (x[52]);
  assign t[632] = (x[31]);
  assign t[633] = (x[32]);
  assign t[634] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[635] = (x[60]);
  assign t[636] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[637] = (x[68]);
  assign t[638] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[639] = (x[74]);
  assign t[63] = ~(t[99] ^ t[100]);
  assign t[640] = (x[23]);
  assign t[641] = (x[39]);
  assign t[642] = (x[40]);
  assign t[643] = (x[47]);
  assign t[644] = (x[48]);
  assign t[645] = (x[53]);
  assign t[646] = (x[54]);
  assign t[647] = (x[88] & ~x[89] & ~x[90] & ~x[91]) | (~x[88] & x[89] & ~x[90] & ~x[91]) | (~x[88] & ~x[89] & x[90] & ~x[91]) | (~x[88] & ~x[89] & ~x[90] & x[91]) | (x[88] & x[89] & x[90] & ~x[91]) | (x[88] & x[89] & ~x[90] & x[91]) | (x[88] & ~x[89] & x[90] & x[91]) | (~x[88] & x[89] & x[90] & x[91]);
  assign t[648] = (x[89]);
  assign t[649] = (x[29]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[650] = (x[61]);
  assign t[651] = (x[62]);
  assign t[652] = (x[69]);
  assign t[653] = (x[70]);
  assign t[654] = (x[101] & ~x[102] & ~x[103] & ~x[104]) | (~x[101] & x[102] & ~x[103] & ~x[104]) | (~x[101] & ~x[102] & x[103] & ~x[104]) | (~x[101] & ~x[102] & ~x[103] & x[104]) | (x[101] & x[102] & x[103] & ~x[104]) | (x[101] & x[102] & ~x[103] & x[104]) | (x[101] & ~x[102] & x[103] & x[104]) | (~x[101] & x[102] & x[103] & x[104]);
  assign t[655] = (x[102]);
  assign t[656] = (x[75]);
  assign t[657] = (x[76]);
  assign t[658] = (x[37]);
  assign t[659] = (x[45]);
  assign t[65] = ~(t[414] | t[103]);
  assign t[660] = (x[51]);
  assign t[661] = (x[90]);
  assign t[662] = (x[91]);
  assign t[663] = (x[59]);
  assign t[664] = (x[67]);
  assign t[665] = (x[103]);
  assign t[666] = (x[104]);
  assign t[667] = (x[73]);
  assign t[668] = (x[88]);
  assign t[669] = (x[101]);
  assign t[66] = ~(t[104] | t[105]);
  assign t[670] = (x[1]);
  assign t[671] = (x[2]);
  assign t[672] = (x[3]);
  assign t[67] = ~(t[106] ^ t[107]);
  assign t[68] = ~(t[415]);
  assign t[69] = ~(t[416]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[110] | t[111]);
  assign t[72] = ~(t[417] | t[112]);
  assign t[73] = t[30] ? x[66] : x[65];
  assign t[74] = ~(t[82] & t[113]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[418] | t[116]);
  assign t[77] = ~(t[117] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[419] | t[123]);
  assign t[81] = ~(t[124] ^ t[125]);
  assign t[82] = ~(t[126] | t[127]);
  assign t[83] = ~(t[128] & t[129]);
  assign t[84] = ~(t[130] & t[131]);
  assign t[85] = t[128] | t[132];
  assign t[86] = ~(t[128]);
  assign t[87] = t[404] ? t[134] : t[133];
  assign t[88] = t[404] ? t[136] : t[135];
  assign t[89] = ~(t[420]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[410] | t[411]);
  assign t[91] = ~(t[421]);
  assign t[92] = ~(t[422]);
  assign t[93] = ~(t[137] | t[138]);
  assign t[94] = ~(t[52] | t[50]);
  assign t[95] = ~(t[139] & t[140]);
  assign t[96] = ~(t[423]);
  assign t[97] = ~(t[424]);
  assign t[98] = ~(t[141] | t[142]);
  assign t[99] = t[143] ? x[85] : x[84];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[205] & ~t[275] & ~t[354]) | (~t[0] & t[205] & ~t[275] & ~t[354]) | (~t[0] & ~t[205] & t[275] & ~t[354]) | (~t[0] & ~t[205] & ~t[275] & t[354]) | (t[0] & t[205] & t[275] & ~t[354]) | (t[0] & t[205] & ~t[275] & t[354]) | (t[0] & ~t[205] & t[275] & t[354]) | (~t[0] & t[205] & t[275] & t[354]);
endmodule

module R2ind131(x, y);
 input [124:0] x;
 output y;

 wire [364:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[108] | t[99]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[109] | t[104]);
  assign t[107] = ~(t[152]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[5];
  assign t[156] = t[201] ^ x[13];
  assign t[157] = t[202] ^ x[16];
  assign t[158] = t[203] ^ x[19];
  assign t[159] = t[204] ^ x[22];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[28];
  assign t[161] = t[206] ^ x[36];
  assign t[162] = t[207] ^ x[39];
  assign t[163] = t[208] ^ x[40];
  assign t[164] = t[209] ^ x[46];
  assign t[165] = t[210] ^ x[52];
  assign t[166] = t[211] ^ x[60];
  assign t[167] = t[212] ^ x[63];
  assign t[168] = t[213] ^ x[64];
  assign t[169] = t[214] ^ x[70];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[76];
  assign t[171] = t[216] ^ x[84];
  assign t[172] = t[217] ^ x[87];
  assign t[173] = t[218] ^ x[88];
  assign t[174] = t[219] ^ x[89];
  assign t[175] = t[220] ^ x[90];
  assign t[176] = t[221] ^ x[91];
  assign t[177] = t[222] ^ x[92];
  assign t[178] = t[223] ^ x[93];
  assign t[179] = t[224] ^ x[99];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[100];
  assign t[181] = t[226] ^ x[101];
  assign t[182] = t[227] ^ x[102];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[104];
  assign t[185] = t[230] ^ x[110];
  assign t[186] = t[231] ^ x[111];
  assign t[187] = t[232] ^ x[112];
  assign t[188] = t[233] ^ x[113];
  assign t[189] = t[234] ^ x[114];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[115];
  assign t[191] = t[236] ^ x[116];
  assign t[192] = t[237] ^ x[117];
  assign t[193] = t[238] ^ x[118];
  assign t[194] = t[239] ^ x[119];
  assign t[195] = t[240] ^ x[120];
  assign t[196] = t[241] ^ x[121];
  assign t[197] = t[242] ^ x[122];
  assign t[198] = t[243] ^ x[123];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[245] & t[246]);
  assign t[201] = (~t[247] & t[248]);
  assign t[202] = (~t[249] & t[250]);
  assign t[203] = (~t[251] & t[252]);
  assign t[204] = (~t[253] & t[254]);
  assign t[205] = (~t[255] & t[256]);
  assign t[206] = (~t[257] & t[258]);
  assign t[207] = (~t[255] & t[259]);
  assign t[208] = (~t[255] & t[260]);
  assign t[209] = (~t[261] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[263] & t[264]);
  assign t[211] = (~t[265] & t[266]);
  assign t[212] = (~t[257] & t[267]);
  assign t[213] = (~t[257] & t[268]);
  assign t[214] = (~t[269] & t[270]);
  assign t[215] = (~t[271] & t[272]);
  assign t[216] = (~t[273] & t[274]);
  assign t[217] = (~t[255] & t[275]);
  assign t[218] = (~t[261] & t[276]);
  assign t[219] = (~t[261] & t[277]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[263] & t[278]);
  assign t[221] = (~t[263] & t[279]);
  assign t[222] = (~t[265] & t[280]);
  assign t[223] = (~t[265] & t[281]);
  assign t[224] = (~t[282] & t[283]);
  assign t[225] = (~t[257] & t[284]);
  assign t[226] = (~t[269] & t[285]);
  assign t[227] = (~t[269] & t[286]);
  assign t[228] = (~t[271] & t[287]);
  assign t[229] = (~t[271] & t[288]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[289] & t[290]);
  assign t[231] = (~t[273] & t[291]);
  assign t[232] = (~t[273] & t[292]);
  assign t[233] = (~t[261] & t[293]);
  assign t[234] = (~t[263] & t[294]);
  assign t[235] = (~t[265] & t[295]);
  assign t[236] = (~t[282] & t[296]);
  assign t[237] = (~t[282] & t[297]);
  assign t[238] = (~t[269] & t[298]);
  assign t[239] = (~t[271] & t[299]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[289] & t[300]);
  assign t[241] = (~t[289] & t[301]);
  assign t[242] = (~t[273] & t[302]);
  assign t[243] = (~t[282] & t[303]);
  assign t[244] = (~t[289] & t[304]);
  assign t[245] = t[305] ^ x[4];
  assign t[246] = t[306] ^ x[5];
  assign t[247] = t[307] ^ x[12];
  assign t[248] = t[308] ^ x[13];
  assign t[249] = t[309] ^ x[15];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[310] ^ x[16];
  assign t[251] = t[311] ^ x[18];
  assign t[252] = t[312] ^ x[19];
  assign t[253] = t[313] ^ x[21];
  assign t[254] = t[314] ^ x[22];
  assign t[255] = t[315] ^ x[27];
  assign t[256] = t[316] ^ x[28];
  assign t[257] = t[317] ^ x[35];
  assign t[258] = t[318] ^ x[36];
  assign t[259] = t[319] ^ x[39];
  assign t[25] = ~(t[113]);
  assign t[260] = t[320] ^ x[40];
  assign t[261] = t[321] ^ x[45];
  assign t[262] = t[322] ^ x[46];
  assign t[263] = t[323] ^ x[51];
  assign t[264] = t[324] ^ x[52];
  assign t[265] = t[325] ^ x[59];
  assign t[266] = t[326] ^ x[60];
  assign t[267] = t[327] ^ x[63];
  assign t[268] = t[328] ^ x[64];
  assign t[269] = t[329] ^ x[69];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[70];
  assign t[271] = t[331] ^ x[75];
  assign t[272] = t[332] ^ x[76];
  assign t[273] = t[333] ^ x[83];
  assign t[274] = t[334] ^ x[84];
  assign t[275] = t[335] ^ x[87];
  assign t[276] = t[336] ^ x[88];
  assign t[277] = t[337] ^ x[89];
  assign t[278] = t[338] ^ x[90];
  assign t[279] = t[339] ^ x[91];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[92];
  assign t[281] = t[341] ^ x[93];
  assign t[282] = t[342] ^ x[98];
  assign t[283] = t[343] ^ x[99];
  assign t[284] = t[344] ^ x[100];
  assign t[285] = t[345] ^ x[101];
  assign t[286] = t[346] ^ x[102];
  assign t[287] = t[347] ^ x[103];
  assign t[288] = t[348] ^ x[104];
  assign t[289] = t[349] ^ x[109];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[110];
  assign t[291] = t[351] ^ x[111];
  assign t[292] = t[352] ^ x[112];
  assign t[293] = t[353] ^ x[113];
  assign t[294] = t[354] ^ x[114];
  assign t[295] = t[355] ^ x[115];
  assign t[296] = t[356] ^ x[116];
  assign t[297] = t[357] ^ x[117];
  assign t[298] = t[358] ^ x[118];
  assign t[299] = t[359] ^ x[119];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[120];
  assign t[301] = t[361] ^ x[121];
  assign t[302] = t[362] ^ x[122];
  assign t[303] = t[363] ^ x[123];
  assign t[304] = t[364] ^ x[124];
  assign t[305] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[306] = (x[3]);
  assign t[307] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[308] = (x[11]);
  assign t[309] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = (x[14]);
  assign t[311] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[312] = (x[17]);
  assign t[313] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[314] = (x[20]);
  assign t[315] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[316] = (x[24]);
  assign t[317] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[318] = (x[32]);
  assign t[319] = (x[26]);
  assign t[31] = t[48] | t[115];
  assign t[320] = (x[23]);
  assign t[321] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[322] = (x[42]);
  assign t[323] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[324] = (x[48]);
  assign t[325] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[326] = (x[56]);
  assign t[327] = (x[34]);
  assign t[328] = (x[31]);
  assign t[329] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[32] = t[18] ? x[30] : x[29];
  assign t[330] = (x[66]);
  assign t[331] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[332] = (x[72]);
  assign t[333] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[334] = (x[80]);
  assign t[335] = (x[25]);
  assign t[336] = (x[44]);
  assign t[337] = (x[41]);
  assign t[338] = (x[50]);
  assign t[339] = (x[47]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[58]);
  assign t[341] = (x[55]);
  assign t[342] = (x[94] & ~x[95] & ~x[96] & ~x[97]) | (~x[94] & x[95] & ~x[96] & ~x[97]) | (~x[94] & ~x[95] & x[96] & ~x[97]) | (~x[94] & ~x[95] & ~x[96] & x[97]) | (x[94] & x[95] & x[96] & ~x[97]) | (x[94] & x[95] & ~x[96] & x[97]) | (x[94] & ~x[95] & x[96] & x[97]) | (~x[94] & x[95] & x[96] & x[97]);
  assign t[343] = (x[95]);
  assign t[344] = (x[33]);
  assign t[345] = (x[68]);
  assign t[346] = (x[65]);
  assign t[347] = (x[74]);
  assign t[348] = (x[71]);
  assign t[349] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[106]);
  assign t[351] = (x[82]);
  assign t[352] = (x[79]);
  assign t[353] = (x[43]);
  assign t[354] = (x[49]);
  assign t[355] = (x[57]);
  assign t[356] = (x[97]);
  assign t[357] = (x[94]);
  assign t[358] = (x[67]);
  assign t[359] = (x[73]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[108]);
  assign t[361] = (x[105]);
  assign t[362] = (x[81]);
  assign t[363] = (x[96]);
  assign t[364] = (x[107]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[57];
  assign t[38] = ~(t[58] & t[59]);
  assign t[39] = t[60] | t[116];
  assign t[3] = ~(t[6]);
  assign t[40] = t[61] ? x[38] : x[37];
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[42];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[74] | t[119];
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = t[77] | t[120];
  assign t[53] = t[78] ? x[54] : x[53];
  assign t[54] = ~(t[79] & t[80]);
  assign t[55] = t[81] | t[121];
  assign t[56] = t[78] ? x[62] : x[61];
  assign t[57] = ~(t[82] & t[83]);
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[123]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[84] | t[58]);
  assign t[61] = ~(t[25]);
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = t[87] | t[124];
  assign t[64] = ~(t[88] & t[89]);
  assign t[65] = t[90] | t[125];
  assign t[66] = t[18] ? x[78] : x[77];
  assign t[67] = ~(t[91] & t[92]);
  assign t[68] = ~(t[93] & t[94]);
  assign t[69] = t[95] | t[126];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[18] ? x[86] : x[85];
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[25]);
  assign t[79] = ~(t[132]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[98] | t[79]);
  assign t[82] = ~(t[99] & t[100]);
  assign t[83] = t[101] | t[134];
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[137]);
  assign t[87] = ~(t[102] | t[85]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[139]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[103] | t[88]);
  assign t[91] = ~(t[104] & t[105]);
  assign t[92] = t[106] | t[140];
  assign t[93] = ~(t[141]);
  assign t[94] = ~(t[142]);
  assign t[95] = ~(t[107] | t[93]);
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [124:0] x;
 output y;

 wire [373:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[142] & t[141]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[155]);
  assign t[104] = ~(t[156]);
  assign t[105] = ~(t[115] & t[116]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[159]);
  assign t[111] = ~(t[160]);
  assign t[112] = ~(t[117] & t[118]);
  assign t[113] = ~(t[151] & t[150]);
  assign t[114] = ~(t[161]);
  assign t[115] = ~(t[156] & t[155]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[160] & t[159]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[5];
  assign t[165] = t[210] ^ x[13];
  assign t[166] = t[211] ^ x[16];
  assign t[167] = t[212] ^ x[19];
  assign t[168] = t[213] ^ x[22];
  assign t[169] = t[214] ^ x[28];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[36];
  assign t[171] = t[216] ^ x[39];
  assign t[172] = t[217] ^ x[40];
  assign t[173] = t[218] ^ x[46];
  assign t[174] = t[219] ^ x[52];
  assign t[175] = t[220] ^ x[60];
  assign t[176] = t[221] ^ x[63];
  assign t[177] = t[222] ^ x[64];
  assign t[178] = t[223] ^ x[70];
  assign t[179] = t[224] ^ x[76];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[84];
  assign t[181] = t[226] ^ x[87];
  assign t[182] = t[227] ^ x[88];
  assign t[183] = t[228] ^ x[89];
  assign t[184] = t[229] ^ x[90];
  assign t[185] = t[230] ^ x[91];
  assign t[186] = t[231] ^ x[92];
  assign t[187] = t[232] ^ x[93];
  assign t[188] = t[233] ^ x[99];
  assign t[189] = t[234] ^ x[100];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[101];
  assign t[191] = t[236] ^ x[102];
  assign t[192] = t[237] ^ x[103];
  assign t[193] = t[238] ^ x[104];
  assign t[194] = t[239] ^ x[110];
  assign t[195] = t[240] ^ x[111];
  assign t[196] = t[241] ^ x[112];
  assign t[197] = t[242] ^ x[113];
  assign t[198] = t[243] ^ x[114];
  assign t[199] = t[244] ^ x[115];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[116];
  assign t[201] = t[246] ^ x[117];
  assign t[202] = t[247] ^ x[118];
  assign t[203] = t[248] ^ x[119];
  assign t[204] = t[249] ^ x[120];
  assign t[205] = t[250] ^ x[121];
  assign t[206] = t[251] ^ x[122];
  assign t[207] = t[252] ^ x[123];
  assign t[208] = t[253] ^ x[124];
  assign t[209] = (~t[254] & t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[256] & t[257]);
  assign t[211] = (~t[258] & t[259]);
  assign t[212] = (~t[260] & t[261]);
  assign t[213] = (~t[262] & t[263]);
  assign t[214] = (~t[264] & t[265]);
  assign t[215] = (~t[266] & t[267]);
  assign t[216] = (~t[264] & t[268]);
  assign t[217] = (~t[264] & t[269]);
  assign t[218] = (~t[270] & t[271]);
  assign t[219] = (~t[272] & t[273]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[274] & t[275]);
  assign t[221] = (~t[266] & t[276]);
  assign t[222] = (~t[266] & t[277]);
  assign t[223] = (~t[278] & t[279]);
  assign t[224] = (~t[280] & t[281]);
  assign t[225] = (~t[282] & t[283]);
  assign t[226] = (~t[264] & t[284]);
  assign t[227] = (~t[270] & t[285]);
  assign t[228] = (~t[270] & t[286]);
  assign t[229] = (~t[272] & t[287]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[272] & t[288]);
  assign t[231] = (~t[274] & t[289]);
  assign t[232] = (~t[274] & t[290]);
  assign t[233] = (~t[291] & t[292]);
  assign t[234] = (~t[266] & t[293]);
  assign t[235] = (~t[278] & t[294]);
  assign t[236] = (~t[278] & t[295]);
  assign t[237] = (~t[280] & t[296]);
  assign t[238] = (~t[280] & t[297]);
  assign t[239] = (~t[298] & t[299]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[282] & t[300]);
  assign t[241] = (~t[282] & t[301]);
  assign t[242] = (~t[270] & t[302]);
  assign t[243] = (~t[272] & t[303]);
  assign t[244] = (~t[274] & t[304]);
  assign t[245] = (~t[291] & t[305]);
  assign t[246] = (~t[291] & t[306]);
  assign t[247] = (~t[278] & t[307]);
  assign t[248] = (~t[280] & t[308]);
  assign t[249] = (~t[298] & t[309]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = (~t[298] & t[310]);
  assign t[251] = (~t[282] & t[311]);
  assign t[252] = (~t[291] & t[312]);
  assign t[253] = (~t[298] & t[313]);
  assign t[254] = t[314] ^ x[4];
  assign t[255] = t[315] ^ x[5];
  assign t[256] = t[316] ^ x[12];
  assign t[257] = t[317] ^ x[13];
  assign t[258] = t[318] ^ x[15];
  assign t[259] = t[319] ^ x[16];
  assign t[25] = ~(t[122]);
  assign t[260] = t[320] ^ x[18];
  assign t[261] = t[321] ^ x[19];
  assign t[262] = t[322] ^ x[21];
  assign t[263] = t[323] ^ x[22];
  assign t[264] = t[324] ^ x[27];
  assign t[265] = t[325] ^ x[28];
  assign t[266] = t[326] ^ x[35];
  assign t[267] = t[327] ^ x[36];
  assign t[268] = t[328] ^ x[39];
  assign t[269] = t[329] ^ x[40];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[45];
  assign t[271] = t[331] ^ x[46];
  assign t[272] = t[332] ^ x[51];
  assign t[273] = t[333] ^ x[52];
  assign t[274] = t[334] ^ x[59];
  assign t[275] = t[335] ^ x[60];
  assign t[276] = t[336] ^ x[63];
  assign t[277] = t[337] ^ x[64];
  assign t[278] = t[338] ^ x[69];
  assign t[279] = t[339] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[75];
  assign t[281] = t[341] ^ x[76];
  assign t[282] = t[342] ^ x[83];
  assign t[283] = t[343] ^ x[84];
  assign t[284] = t[344] ^ x[87];
  assign t[285] = t[345] ^ x[88];
  assign t[286] = t[346] ^ x[89];
  assign t[287] = t[347] ^ x[90];
  assign t[288] = t[348] ^ x[91];
  assign t[289] = t[349] ^ x[92];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[93];
  assign t[291] = t[351] ^ x[98];
  assign t[292] = t[352] ^ x[99];
  assign t[293] = t[353] ^ x[100];
  assign t[294] = t[354] ^ x[101];
  assign t[295] = t[355] ^ x[102];
  assign t[296] = t[356] ^ x[103];
  assign t[297] = t[357] ^ x[104];
  assign t[298] = t[358] ^ x[109];
  assign t[299] = t[359] ^ x[110];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[111];
  assign t[301] = t[361] ^ x[112];
  assign t[302] = t[362] ^ x[113];
  assign t[303] = t[363] ^ x[114];
  assign t[304] = t[364] ^ x[115];
  assign t[305] = t[365] ^ x[116];
  assign t[306] = t[366] ^ x[117];
  assign t[307] = t[367] ^ x[118];
  assign t[308] = t[368] ^ x[119];
  assign t[309] = t[369] ^ x[120];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[370] ^ x[121];
  assign t[311] = t[371] ^ x[122];
  assign t[312] = t[372] ^ x[123];
  assign t[313] = t[373] ^ x[124];
  assign t[314] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[315] = (x[2]);
  assign t[316] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[317] = (x[11]);
  assign t[318] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[319] = (x[14]);
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[321] = (x[17]);
  assign t[322] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[323] = (x[20]);
  assign t[324] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[325] = (x[24]);
  assign t[326] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[327] = (x[32]);
  assign t[328] = (x[26]);
  assign t[329] = (x[23]);
  assign t[32] = t[18] ? x[30] : x[29];
  assign t[330] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[331] = (x[42]);
  assign t[332] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[333] = (x[48]);
  assign t[334] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[335] = (x[56]);
  assign t[336] = (x[34]);
  assign t[337] = (x[31]);
  assign t[338] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[339] = (x[66]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[341] = (x[72]);
  assign t[342] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[343] = (x[80]);
  assign t[344] = (x[25]);
  assign t[345] = (x[44]);
  assign t[346] = (x[41]);
  assign t[347] = (x[50]);
  assign t[348] = (x[47]);
  assign t[349] = (x[58]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[55]);
  assign t[351] = (x[94] & ~x[95] & ~x[96] & ~x[97]) | (~x[94] & x[95] & ~x[96] & ~x[97]) | (~x[94] & ~x[95] & x[96] & ~x[97]) | (~x[94] & ~x[95] & ~x[96] & x[97]) | (x[94] & x[95] & x[96] & ~x[97]) | (x[94] & x[95] & ~x[96] & x[97]) | (x[94] & ~x[95] & x[96] & x[97]) | (~x[94] & x[95] & x[96] & x[97]);
  assign t[352] = (x[95]);
  assign t[353] = (x[33]);
  assign t[354] = (x[68]);
  assign t[355] = (x[65]);
  assign t[356] = (x[74]);
  assign t[357] = (x[71]);
  assign t[358] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[359] = (x[106]);
  assign t[35] = t[53] ^ t[36];
  assign t[360] = (x[82]);
  assign t[361] = (x[79]);
  assign t[362] = (x[43]);
  assign t[363] = (x[49]);
  assign t[364] = (x[57]);
  assign t[365] = (x[97]);
  assign t[366] = (x[94]);
  assign t[367] = (x[67]);
  assign t[368] = (x[73]);
  assign t[369] = (x[108]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[105]);
  assign t[371] = (x[81]);
  assign t[372] = (x[96]);
  assign t[373] = (x[107]);
  assign t[37] = t[56] ^ t[57];
  assign t[38] = ~(t[58] & t[59]);
  assign t[39] = ~(t[60] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[61] ? x[38] : x[37];
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[42];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[75] & t[128]);
  assign t[51] = ~(t[76] & t[77]);
  assign t[52] = ~(t[78] & t[129]);
  assign t[53] = t[61] ? x[54] : x[53];
  assign t[54] = ~(t[79] & t[80]);
  assign t[55] = ~(t[81] & t[130]);
  assign t[56] = t[61] ? x[62] : x[61];
  assign t[57] = ~(t[82] & t[83]);
  assign t[58] = ~(t[131]);
  assign t[59] = ~(t[132]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[84] & t[85]);
  assign t[61] = ~(t[25]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[133]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[134]);
  assign t[66] = t[18] ? x[78] : x[77];
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = ~(t[94] & t[95]);
  assign t[69] = ~(t[96] & t[135]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[122] ? x[86] : x[85];
  assign t[71] = ~(t[127] & t[126]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[97] & t[98]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[141]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[142]);
  assign t[81] = ~(t[101] & t[102]);
  assign t[82] = ~(t[103] & t[104]);
  assign t[83] = ~(t[105] & t[143]);
  assign t[84] = ~(t[132] & t[131]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[147]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[108] & t[109]);
  assign t[92] = ~(t[110] & t[111]);
  assign t[93] = ~(t[112] & t[149]);
  assign t[94] = ~(t[150]);
  assign t[95] = ~(t[151]);
  assign t[96] = ~(t[113] & t[114]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [114:0] x;
 output y;

 wire [304:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[5];
  assign t[136] = t[171] ^ x[13];
  assign t[137] = t[172] ^ x[16];
  assign t[138] = t[173] ^ x[19];
  assign t[139] = t[174] ^ x[22];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[28];
  assign t[141] = t[176] ^ x[29];
  assign t[142] = t[177] ^ x[37];
  assign t[143] = t[178] ^ x[38];
  assign t[144] = t[179] ^ x[41];
  assign t[145] = t[180] ^ x[47];
  assign t[146] = t[181] ^ x[48];
  assign t[147] = t[182] ^ x[54];
  assign t[148] = t[183] ^ x[55];
  assign t[149] = t[184] ^ x[63];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[64];
  assign t[151] = t[186] ^ x[67];
  assign t[152] = t[187] ^ x[73];
  assign t[153] = t[188] ^ x[74];
  assign t[154] = t[189] ^ x[80];
  assign t[155] = t[190] ^ x[81];
  assign t[156] = t[191] ^ x[89];
  assign t[157] = t[192] ^ x[90];
  assign t[158] = t[193] ^ x[93];
  assign t[159] = t[194] ^ x[94];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[100];
  assign t[161] = t[196] ^ x[101];
  assign t[162] = t[197] ^ x[102];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[104];
  assign t[165] = t[200] ^ x[105];
  assign t[166] = t[201] ^ x[111];
  assign t[167] = t[202] ^ x[112];
  assign t[168] = t[203] ^ x[113];
  assign t[169] = t[204] ^ x[114];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (~t[205] & t[206]);
  assign t[171] = (~t[207] & t[208]);
  assign t[172] = (~t[209] & t[210]);
  assign t[173] = (~t[211] & t[212]);
  assign t[174] = (~t[213] & t[214]);
  assign t[175] = (~t[215] & t[216]);
  assign t[176] = (~t[215] & t[217]);
  assign t[177] = (~t[218] & t[219]);
  assign t[178] = (~t[218] & t[220]);
  assign t[179] = (~t[215] & t[221]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (~t[222] & t[223]);
  assign t[181] = (~t[222] & t[224]);
  assign t[182] = (~t[225] & t[226]);
  assign t[183] = (~t[225] & t[227]);
  assign t[184] = (~t[228] & t[229]);
  assign t[185] = (~t[228] & t[230]);
  assign t[186] = (~t[218] & t[231]);
  assign t[187] = (~t[232] & t[233]);
  assign t[188] = (~t[232] & t[234]);
  assign t[189] = (~t[235] & t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (~t[235] & t[237]);
  assign t[191] = (~t[238] & t[239]);
  assign t[192] = (~t[238] & t[240]);
  assign t[193] = (~t[222] & t[241]);
  assign t[194] = (~t[225] & t[242]);
  assign t[195] = (~t[243] & t[244]);
  assign t[196] = (~t[243] & t[245]);
  assign t[197] = (~t[228] & t[246]);
  assign t[198] = (~t[232] & t[247]);
  assign t[199] = (~t[235] & t[248]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[238] & t[249]);
  assign t[201] = (~t[250] & t[251]);
  assign t[202] = (~t[250] & t[252]);
  assign t[203] = (~t[243] & t[253]);
  assign t[204] = (~t[250] & t[254]);
  assign t[205] = t[255] ^ x[4];
  assign t[206] = t[256] ^ x[5];
  assign t[207] = t[257] ^ x[12];
  assign t[208] = t[258] ^ x[13];
  assign t[209] = t[259] ^ x[15];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[260] ^ x[16];
  assign t[211] = t[261] ^ x[18];
  assign t[212] = t[262] ^ x[19];
  assign t[213] = t[263] ^ x[21];
  assign t[214] = t[264] ^ x[22];
  assign t[215] = t[265] ^ x[27];
  assign t[216] = t[266] ^ x[28];
  assign t[217] = t[267] ^ x[29];
  assign t[218] = t[268] ^ x[36];
  assign t[219] = t[269] ^ x[37];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[270] ^ x[38];
  assign t[221] = t[271] ^ x[41];
  assign t[222] = t[272] ^ x[46];
  assign t[223] = t[273] ^ x[47];
  assign t[224] = t[274] ^ x[48];
  assign t[225] = t[275] ^ x[53];
  assign t[226] = t[276] ^ x[54];
  assign t[227] = t[277] ^ x[55];
  assign t[228] = t[278] ^ x[62];
  assign t[229] = t[279] ^ x[63];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[280] ^ x[64];
  assign t[231] = t[281] ^ x[67];
  assign t[232] = t[282] ^ x[72];
  assign t[233] = t[283] ^ x[73];
  assign t[234] = t[284] ^ x[74];
  assign t[235] = t[285] ^ x[79];
  assign t[236] = t[286] ^ x[80];
  assign t[237] = t[287] ^ x[81];
  assign t[238] = t[288] ^ x[88];
  assign t[239] = t[289] ^ x[89];
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = t[290] ^ x[90];
  assign t[241] = t[291] ^ x[93];
  assign t[242] = t[292] ^ x[94];
  assign t[243] = t[293] ^ x[99];
  assign t[244] = t[294] ^ x[100];
  assign t[245] = t[295] ^ x[101];
  assign t[246] = t[296] ^ x[102];
  assign t[247] = t[297] ^ x[103];
  assign t[248] = t[298] ^ x[104];
  assign t[249] = t[299] ^ x[105];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[300] ^ x[110];
  assign t[251] = t[301] ^ x[111];
  assign t[252] = t[302] ^ x[112];
  assign t[253] = t[303] ^ x[113];
  assign t[254] = t[304] ^ x[114];
  assign t[255] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[256] = (x[1]);
  assign t[257] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[258] = (x[11]);
  assign t[259] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[25] = ~(t[103]);
  assign t[260] = (x[14]);
  assign t[261] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[262] = (x[17]);
  assign t[263] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[264] = (x[20]);
  assign t[265] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[266] = (x[25]);
  assign t[267] = (x[23]);
  assign t[268] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[269] = (x[34]);
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = (x[32]);
  assign t[271] = (x[26]);
  assign t[272] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[273] = (x[44]);
  assign t[274] = (x[42]);
  assign t[275] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[276] = (x[51]);
  assign t[277] = (x[49]);
  assign t[278] = (x[58] & ~x[59] & ~x[60] & ~x[61]) | (~x[58] & x[59] & ~x[60] & ~x[61]) | (~x[58] & ~x[59] & x[60] & ~x[61]) | (~x[58] & ~x[59] & ~x[60] & x[61]) | (x[58] & x[59] & x[60] & ~x[61]) | (x[58] & x[59] & ~x[60] & x[61]) | (x[58] & ~x[59] & x[60] & x[61]) | (~x[58] & x[59] & x[60] & x[61]);
  assign t[279] = (x[60]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[58]);
  assign t[281] = (x[35]);
  assign t[282] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[283] = (x[70]);
  assign t[284] = (x[68]);
  assign t[285] = (x[75] & ~x[76] & ~x[77] & ~x[78]) | (~x[75] & x[76] & ~x[77] & ~x[78]) | (~x[75] & ~x[76] & x[77] & ~x[78]) | (~x[75] & ~x[76] & ~x[77] & x[78]) | (x[75] & x[76] & x[77] & ~x[78]) | (x[75] & x[76] & ~x[77] & x[78]) | (x[75] & ~x[76] & x[77] & x[78]) | (~x[75] & x[76] & x[77] & x[78]);
  assign t[286] = (x[77]);
  assign t[287] = (x[75]);
  assign t[288] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[289] = (x[86]);
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = (x[84]);
  assign t[291] = (x[45]);
  assign t[292] = (x[52]);
  assign t[293] = (x[95] & ~x[96] & ~x[97] & ~x[98]) | (~x[95] & x[96] & ~x[97] & ~x[98]) | (~x[95] & ~x[96] & x[97] & ~x[98]) | (~x[95] & ~x[96] & ~x[97] & x[98]) | (x[95] & x[96] & x[97] & ~x[98]) | (x[95] & x[96] & ~x[97] & x[98]) | (x[95] & ~x[96] & x[97] & x[98]) | (~x[95] & x[96] & x[97] & x[98]);
  assign t[294] = (x[97]);
  assign t[295] = (x[95]);
  assign t[296] = (x[61]);
  assign t[297] = (x[71]);
  assign t[298] = (x[78]);
  assign t[299] = (x[87]);
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[106] & ~x[107] & ~x[108] & ~x[109]) | (~x[106] & x[107] & ~x[108] & ~x[109]) | (~x[106] & ~x[107] & x[108] & ~x[109]) | (~x[106] & ~x[107] & ~x[108] & x[109]) | (x[106] & x[107] & x[108] & ~x[109]) | (x[106] & x[107] & ~x[108] & x[109]) | (x[106] & ~x[107] & x[108] & x[109]) | (~x[106] & x[107] & x[108] & x[109]);
  assign t[301] = (x[108]);
  assign t[302] = (x[106]);
  assign t[303] = (x[98]);
  assign t[304] = (x[109]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[32] = t[48] ? x[31] : x[30];
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[54];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[34];
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = ~(t[108] & t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[48] ? x[40] : x[39];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[44];
  assign t[44] = ~(t[65] & t[66]);
  assign t[45] = t[67] ^ t[68];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[69]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = ~(t[113] & t[73]);
  assign t[53] = t[74] ? x[57] : x[56];
  assign t[54] = ~(t[75] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = ~(t[115] & t[78]);
  assign t[57] = t[74] ? x[66] : x[65];
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = ~(t[120] & t[83]);
  assign t[64] = t[74] ? x[83] : x[82];
  assign t[65] = ~(t[121] & t[84]);
  assign t[66] = ~(t[122] & t[85]);
  assign t[67] = t[48] ? x[92] : x[91];
  assign t[68] = ~(t[86] & t[87]);
  assign t[69] = ~(t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[123]);
  assign t[71] = ~(t[123] & t[88]);
  assign t[72] = ~(t[124]);
  assign t[73] = ~(t[124] & t[89]);
  assign t[74] = ~(t[25]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126] & t[91]);
  assign t[77] = ~(t[127]);
  assign t[78] = ~(t[127] & t[92]);
  assign t[79] = ~(t[107]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[128]);
  assign t[81] = ~(t[128] & t[93]);
  assign t[82] = ~(t[129]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[133] & t[98]);
  assign t[92] = ~(t[114]);
  assign t[93] = ~(t[117]);
  assign t[94] = ~(t[119]);
  assign t[95] = ~(t[121]);
  assign t[96] = ~(t[134]);
  assign t[97] = ~(t[134] & t[99]);
  assign t[98] = ~(t[125]);
  assign t[99] = ~(t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [124:0] x;
 output y;

 wire [459:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = t[144] | t[145];
  assign t[101] = ~(t[227]);
  assign t[102] = ~(t[228]);
  assign t[103] = ~(t[146] | t[147]);
  assign t[104] = ~(t[148] | t[149]);
  assign t[105] = ~(t[229] | t[150]);
  assign t[106] = t[143] ? x[95] : x[94];
  assign t[107] = ~(t[151] & t[152]);
  assign t[108] = ~(t[230]);
  assign t[109] = ~(t[217] | t[218]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[232]);
  assign t[112] = ~(t[153] | t[154]);
  assign t[113] = ~(t[155] | t[156]);
  assign t[114] = ~(t[233]);
  assign t[115] = ~(t[234]);
  assign t[116] = ~(t[157] | t[158]);
  assign t[117] = ~(t[159] | t[160]);
  assign t[118] = ~(t[235] | t[161]);
  assign t[119] = t[30] ? x[108] : x[107];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[162] & t[163]);
  assign t[121] = ~(t[236]);
  assign t[122] = ~(t[237]);
  assign t[123] = ~(t[164] | t[165]);
  assign t[124] = t[30] ? x[112] : x[111];
  assign t[125] = ~(t[166] & t[167]);
  assign t[126] = ~(t[128] | t[168]);
  assign t[127] = ~(t[86] | t[169]);
  assign t[128] = ~(t[208]);
  assign t[129] = ~(t[170] & t[171]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[209] & t[172];
  assign t[131] = t[173] | t[174];
  assign t[132] = t[206] ? t[170] : t[175];
  assign t[133] = ~(t[173] & t[176]);
  assign t[134] = ~(t[174] & t[209]);
  assign t[135] = ~(t[173] & t[209]);
  assign t[136] = ~(t[174] & t[176]);
  assign t[137] = ~(t[238]);
  assign t[138] = ~(t[223] | t[224]);
  assign t[139] = ~(t[207] | t[176]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[86] & t[206];
  assign t[141] = ~(t[239]);
  assign t[142] = ~(t[225] | t[226]);
  assign t[143] = ~(t[49]);
  assign t[144] = ~(t[177] & t[95]);
  assign t[145] = ~(t[86] | t[178]);
  assign t[146] = ~(t[240]);
  assign t[147] = ~(t[227] | t[228]);
  assign t[148] = ~(t[241]);
  assign t[149] = ~(t[242]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[179] | t[180]);
  assign t[151] = ~(t[52]);
  assign t[152] = ~(t[181] | t[145]);
  assign t[153] = ~(t[243]);
  assign t[154] = ~(t[231] | t[232]);
  assign t[155] = ~(t[86] | t[182]);
  assign t[156] = ~(t[32] & t[85]);
  assign t[157] = ~(t[244]);
  assign t[158] = ~(t[233] | t[234]);
  assign t[159] = ~(t[245]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[246]);
  assign t[161] = ~(t[183] | t[184]);
  assign t[162] = ~(t[52] | t[185]);
  assign t[163] = ~(t[100] | t[186]);
  assign t[164] = ~(t[247]);
  assign t[165] = ~(t[236] | t[237]);
  assign t[166] = ~(t[187] | t[155]);
  assign t[167] = ~(t[126] | t[144]);
  assign t[168] = t[206] ? t[133] : t[136];
  assign t[169] = t[206] ? t[175] : t[188];
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = ~(x[7] & t[189]);
  assign t[171] = ~(t[209] & t[190]);
  assign t[172] = ~(t[128] | t[206]);
  assign t[173] = ~(x[7] | t[207]);
  assign t[174] = x[7] & t[207];
  assign t[175] = ~(t[190] & t[176]);
  assign t[176] = ~(t[209]);
  assign t[177] = ~(t[191] | t[192]);
  assign t[178] = t[206] ? t[171] : t[170];
  assign t[179] = ~(t[248]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[241] | t[242]);
  assign t[181] = ~(t[193]);
  assign t[182] = t[206] ? t[135] : t[136];
  assign t[183] = ~(t[249]);
  assign t[184] = ~(t[245] | t[246]);
  assign t[185] = ~(t[86] | t[194]);
  assign t[186] = ~(t[195] & t[85]);
  assign t[187] = ~(t[86] | t[196]);
  assign t[188] = ~(x[7] & t[139]);
  assign t[189] = ~(t[207] | t[209]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(x[7] | t[197]);
  assign t[191] = ~(t[128] | t[198]);
  assign t[192] = ~(t[128] | t[199]);
  assign t[193] = ~(t[200] | t[53]);
  assign t[194] = t[206] ? t[170] : t[171];
  assign t[195] = ~(t[201] | t[200]);
  assign t[196] = t[206] ? t[133] : t[134];
  assign t[197] = ~(t[207]);
  assign t[198] = t[206] ? t[136] : t[133];
  assign t[199] = t[206] ? t[175] : t[170];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[86] | t[202]);
  assign t[201] = ~(t[203]);
  assign t[202] = t[206] ? t[188] : t[175];
  assign t[203] = ~(t[172] & t[204]);
  assign t[204] = ~(t[171] & t[188]);
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[9] : x[10];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = t[295] ^ x[5];
  assign t[251] = t[296] ^ x[13];
  assign t[252] = t[297] ^ x[16];
  assign t[253] = t[298] ^ x[19];
  assign t[254] = t[299] ^ x[22];
  assign t[255] = t[300] ^ x[28];
  assign t[256] = t[301] ^ x[34];
  assign t[257] = t[302] ^ x[35];
  assign t[258] = t[303] ^ x[36];
  assign t[259] = t[304] ^ x[42];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[50];
  assign t[261] = t[306] ^ x[56];
  assign t[262] = t[307] ^ x[57];
  assign t[263] = t[308] ^ x[58];
  assign t[264] = t[309] ^ x[64];
  assign t[265] = t[310] ^ x[72];
  assign t[266] = t[311] ^ x[78];
  assign t[267] = t[312] ^ x[79];
  assign t[268] = t[313] ^ x[80];
  assign t[269] = t[314] ^ x[81];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[82];
  assign t[271] = t[316] ^ x[83];
  assign t[272] = t[317] ^ x[86];
  assign t[273] = t[318] ^ x[87];
  assign t[274] = t[319] ^ x[93];
  assign t[275] = t[320] ^ x[96];
  assign t[276] = t[321] ^ x[97];
  assign t[277] = t[322] ^ x[98];
  assign t[278] = t[323] ^ x[99];
  assign t[279] = t[324] ^ x[100];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[106];
  assign t[281] = t[326] ^ x[109];
  assign t[282] = t[327] ^ x[110];
  assign t[283] = t[328] ^ x[113];
  assign t[284] = t[329] ^ x[114];
  assign t[285] = t[330] ^ x[115];
  assign t[286] = t[331] ^ x[116];
  assign t[287] = t[332] ^ x[117];
  assign t[288] = t[333] ^ x[118];
  assign t[289] = t[334] ^ x[119];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[120];
  assign t[291] = t[336] ^ x[121];
  assign t[292] = t[337] ^ x[122];
  assign t[293] = t[338] ^ x[123];
  assign t[294] = t[339] ^ x[124];
  assign t[295] = (~t[340] & t[341]);
  assign t[296] = (~t[342] & t[343]);
  assign t[297] = (~t[344] & t[345]);
  assign t[298] = (~t[346] & t[347]);
  assign t[299] = (~t[348] & t[349]);
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[350] & t[351]);
  assign t[301] = (~t[352] & t[353]);
  assign t[302] = (~t[350] & t[354]);
  assign t[303] = (~t[350] & t[355]);
  assign t[304] = (~t[356] & t[357]);
  assign t[305] = (~t[358] & t[359]);
  assign t[306] = (~t[360] & t[361]);
  assign t[307] = (~t[352] & t[362]);
  assign t[308] = (~t[352] & t[363]);
  assign t[309] = (~t[364] & t[365]);
  assign t[30] = ~(t[49]);
  assign t[310] = (~t[366] & t[367]);
  assign t[311] = (~t[368] & t[369]);
  assign t[312] = (~t[350] & t[370]);
  assign t[313] = (~t[356] & t[371]);
  assign t[314] = (~t[356] & t[372]);
  assign t[315] = (~t[358] & t[373]);
  assign t[316] = (~t[358] & t[374]);
  assign t[317] = (~t[360] & t[375]);
  assign t[318] = (~t[360] & t[376]);
  assign t[319] = (~t[377] & t[378]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (~t[352] & t[379]);
  assign t[321] = (~t[364] & t[380]);
  assign t[322] = (~t[364] & t[381]);
  assign t[323] = (~t[366] & t[382]);
  assign t[324] = (~t[366] & t[383]);
  assign t[325] = (~t[384] & t[385]);
  assign t[326] = (~t[368] & t[386]);
  assign t[327] = (~t[368] & t[387]);
  assign t[328] = (~t[356] & t[388]);
  assign t[329] = (~t[358] & t[389]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (~t[360] & t[390]);
  assign t[331] = (~t[377] & t[391]);
  assign t[332] = (~t[377] & t[392]);
  assign t[333] = (~t[364] & t[393]);
  assign t[334] = (~t[366] & t[394]);
  assign t[335] = (~t[384] & t[395]);
  assign t[336] = (~t[384] & t[396]);
  assign t[337] = (~t[368] & t[397]);
  assign t[338] = (~t[377] & t[398]);
  assign t[339] = (~t[384] & t[399]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = t[400] ^ x[4];
  assign t[341] = t[401] ^ x[5];
  assign t[342] = t[402] ^ x[12];
  assign t[343] = t[403] ^ x[13];
  assign t[344] = t[404] ^ x[15];
  assign t[345] = t[405] ^ x[16];
  assign t[346] = t[406] ^ x[18];
  assign t[347] = t[407] ^ x[19];
  assign t[348] = t[408] ^ x[21];
  assign t[349] = t[409] ^ x[22];
  assign t[34] = ~(t[210] | t[56]);
  assign t[350] = t[410] ^ x[27];
  assign t[351] = t[411] ^ x[28];
  assign t[352] = t[412] ^ x[33];
  assign t[353] = t[413] ^ x[34];
  assign t[354] = t[414] ^ x[35];
  assign t[355] = t[415] ^ x[36];
  assign t[356] = t[416] ^ x[41];
  assign t[357] = t[417] ^ x[42];
  assign t[358] = t[418] ^ x[49];
  assign t[359] = t[419] ^ x[50];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[420] ^ x[55];
  assign t[361] = t[421] ^ x[56];
  assign t[362] = t[422] ^ x[57];
  assign t[363] = t[423] ^ x[58];
  assign t[364] = t[424] ^ x[63];
  assign t[365] = t[425] ^ x[64];
  assign t[366] = t[426] ^ x[71];
  assign t[367] = t[427] ^ x[72];
  assign t[368] = t[428] ^ x[77];
  assign t[369] = t[429] ^ x[78];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[430] ^ x[79];
  assign t[371] = t[431] ^ x[80];
  assign t[372] = t[432] ^ x[81];
  assign t[373] = t[433] ^ x[82];
  assign t[374] = t[434] ^ x[83];
  assign t[375] = t[435] ^ x[86];
  assign t[376] = t[436] ^ x[87];
  assign t[377] = t[437] ^ x[92];
  assign t[378] = t[438] ^ x[93];
  assign t[379] = t[439] ^ x[96];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[440] ^ x[97];
  assign t[381] = t[441] ^ x[98];
  assign t[382] = t[442] ^ x[99];
  assign t[383] = t[443] ^ x[100];
  assign t[384] = t[444] ^ x[105];
  assign t[385] = t[445] ^ x[106];
  assign t[386] = t[446] ^ x[109];
  assign t[387] = t[447] ^ x[110];
  assign t[388] = t[448] ^ x[113];
  assign t[389] = t[449] ^ x[114];
  assign t[38] = ~(t[39] ^ t[63]);
  assign t[390] = t[450] ^ x[115];
  assign t[391] = t[451] ^ x[116];
  assign t[392] = t[452] ^ x[117];
  assign t[393] = t[453] ^ x[118];
  assign t[394] = t[454] ^ x[119];
  assign t[395] = t[455] ^ x[120];
  assign t[396] = t[456] ^ x[121];
  assign t[397] = t[457] ^ x[122];
  assign t[398] = t[458] ^ x[123];
  assign t[399] = t[459] ^ x[124];
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[401] = (x[0]);
  assign t[402] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[403] = (x[11]);
  assign t[404] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[405] = (x[14]);
  assign t[406] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[407] = (x[17]);
  assign t[408] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[409] = (x[20]);
  assign t[40] = ~(t[66] ^ t[67]);
  assign t[410] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[411] = (x[24]);
  assign t[412] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[413] = (x[30]);
  assign t[414] = (x[25]);
  assign t[415] = (x[26]);
  assign t[416] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[417] = (x[38]);
  assign t[418] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[419] = (x[46]);
  assign t[41] = ~(t[68] | t[69]);
  assign t[420] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[421] = (x[52]);
  assign t[422] = (x[31]);
  assign t[423] = (x[32]);
  assign t[424] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[425] = (x[60]);
  assign t[426] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[427] = (x[68]);
  assign t[428] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[429] = (x[74]);
  assign t[42] = ~(t[211] | t[70]);
  assign t[430] = (x[23]);
  assign t[431] = (x[39]);
  assign t[432] = (x[40]);
  assign t[433] = (x[47]);
  assign t[434] = (x[48]);
  assign t[435] = (x[53]);
  assign t[436] = (x[54]);
  assign t[437] = (x[88] & ~x[89] & ~x[90] & ~x[91]) | (~x[88] & x[89] & ~x[90] & ~x[91]) | (~x[88] & ~x[89] & x[90] & ~x[91]) | (~x[88] & ~x[89] & ~x[90] & x[91]) | (x[88] & x[89] & x[90] & ~x[91]) | (x[88] & x[89] & ~x[90] & x[91]) | (x[88] & ~x[89] & x[90] & x[91]) | (~x[88] & x[89] & x[90] & x[91]);
  assign t[438] = (x[89]);
  assign t[439] = (x[29]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[440] = (x[61]);
  assign t[441] = (x[62]);
  assign t[442] = (x[69]);
  assign t[443] = (x[70]);
  assign t[444] = (x[101] & ~x[102] & ~x[103] & ~x[104]) | (~x[101] & x[102] & ~x[103] & ~x[104]) | (~x[101] & ~x[102] & x[103] & ~x[104]) | (~x[101] & ~x[102] & ~x[103] & x[104]) | (x[101] & x[102] & x[103] & ~x[104]) | (x[101] & x[102] & ~x[103] & x[104]) | (x[101] & ~x[102] & x[103] & x[104]) | (~x[101] & x[102] & x[103] & x[104]);
  assign t[445] = (x[102]);
  assign t[446] = (x[75]);
  assign t[447] = (x[76]);
  assign t[448] = (x[37]);
  assign t[449] = (x[45]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[450] = (x[51]);
  assign t[451] = (x[90]);
  assign t[452] = (x[91]);
  assign t[453] = (x[59]);
  assign t[454] = (x[67]);
  assign t[455] = (x[103]);
  assign t[456] = (x[104]);
  assign t[457] = (x[73]);
  assign t[458] = (x[88]);
  assign t[459] = (x[101]);
  assign t[45] = ~(t[75] | t[76]);
  assign t[46] = ~(t[77] ^ t[78]);
  assign t[47] = ~(t[79] | t[80]);
  assign t[48] = ~(t[45] ^ t[81]);
  assign t[49] = ~(t[208]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[82] & t[83]);
  assign t[51] = ~(t[84] & t[85]);
  assign t[52] = ~(t[86] | t[87]);
  assign t[53] = ~(t[86] | t[88]);
  assign t[54] = ~(t[212]);
  assign t[55] = ~(t[213]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[214] | t[93]);
  assign t[59] = t[30] ? x[44] : x[43];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[215] | t[98]);
  assign t[63] = ~(t[99] ^ t[100]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[65] = ~(t[216] | t[103]);
  assign t[66] = ~(t[104] | t[105]);
  assign t[67] = ~(t[106] ^ t[107]);
  assign t[68] = ~(t[217]);
  assign t[69] = ~(t[218]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[110] | t[111]);
  assign t[72] = ~(t[219] | t[112]);
  assign t[73] = t[30] ? x[66] : x[65];
  assign t[74] = ~(t[82] & t[113]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[220] | t[116]);
  assign t[77] = ~(t[117] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[121] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[221] | t[123]);
  assign t[81] = ~(t[124] ^ t[125]);
  assign t[82] = ~(t[126] | t[127]);
  assign t[83] = ~(t[128] & t[129]);
  assign t[84] = ~(t[130] & t[131]);
  assign t[85] = t[128] | t[132];
  assign t[86] = ~(t[128]);
  assign t[87] = t[206] ? t[134] : t[133];
  assign t[88] = t[206] ? t[136] : t[135];
  assign t[89] = ~(t[222]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[212] | t[213]);
  assign t[91] = ~(t[223]);
  assign t[92] = ~(t[224]);
  assign t[93] = ~(t[137] | t[138]);
  assign t[94] = ~(t[52] | t[50]);
  assign t[95] = ~(t[139] & t[140]);
  assign t[96] = ~(t[225]);
  assign t[97] = ~(t[226]);
  assign t[98] = ~(t[141] | t[142]);
  assign t[99] = t[143] ? x[85] : x[84];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [163:0] x;
 output y;

 wire [638:0] t;
  assign t[0] = t[1] ? t[2] : t[391];
  assign t[100] = ~(t[139] | t[140]);
  assign t[101] = t[141] ? x[87] : x[86];
  assign t[102] = ~(t[142] & t[143]);
  assign t[103] = ~(t[413]);
  assign t[104] = ~(t[402] | t[403]);
  assign t[105] = ~(t[414]);
  assign t[106] = ~(t[415]);
  assign t[107] = ~(t[144] | t[145]);
  assign t[108] = ~(t[146] | t[147]);
  assign t[109] = ~(t[416]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[417]);
  assign t[111] = ~(t[148] | t[149]);
  assign t[112] = ~(t[150] | t[151]);
  assign t[113] = ~(t[418] | t[152]);
  assign t[114] = t[30] ? x[100] : x[99];
  assign t[115] = ~(t[153] & t[154]);
  assign t[116] = ~(t[419]);
  assign t[117] = ~(t[420]);
  assign t[118] = ~(t[155] | t[156]);
  assign t[119] = t[30] ? x[104] : x[103];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[157] & t[158]);
  assign t[121] = ~(t[159] & t[160]);
  assign t[122] = ~(t[161] & t[160]);
  assign t[123] = ~(x[7] & t[162]);
  assign t[124] = ~(t[163] & t[160]);
  assign t[125] = ~(t[161] & t[395]);
  assign t[126] = ~(t[81] | t[164]);
  assign t[127] = ~(t[81] | t[165]);
  assign t[128] = t[392] ? t[166] : t[124];
  assign t[129] = ~(t[79] | t[167]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[168]);
  assign t[131] = ~(t[81] | t[169]);
  assign t[132] = ~(t[421]);
  assign t[133] = ~(t[408] | t[409]);
  assign t[134] = ~(t[422]);
  assign t[135] = ~(t[423]);
  assign t[136] = ~(t[170] | t[171]);
  assign t[137] = ~(t[172] | t[127]);
  assign t[138] = ~(t[173] | t[174]);
  assign t[139] = ~(t[424]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[411] | t[412]);
  assign t[141] = ~(t[48]);
  assign t[142] = ~(t[175] | t[176]);
  assign t[143] = ~(t[177]);
  assign t[144] = ~(t[425]);
  assign t[145] = ~(t[414] | t[415]);
  assign t[146] = ~(t[31] & t[178]);
  assign t[147] = ~(t[179] & t[85]);
  assign t[148] = ~(t[426]);
  assign t[149] = ~(t[416] | t[417]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[427]);
  assign t[151] = ~(t[428]);
  assign t[152] = ~(t[180] | t[181]);
  assign t[153] = ~(t[126] | t[172]);
  assign t[154] = ~(t[182] | t[183]);
  assign t[155] = ~(t[429]);
  assign t[156] = ~(t[419] | t[420]);
  assign t[157] = ~(t[177] | t[51]);
  assign t[158] = ~(t[49] | t[184]);
  assign t[159] = x[7] & t[393];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[395]);
  assign t[161] = ~(x[7] | t[393]);
  assign t[162] = ~(t[393] | t[160]);
  assign t[163] = ~(x[7] | t[185]);
  assign t[164] = t[392] ? t[186] : t[122];
  assign t[165] = t[392] ? t[121] : t[125];
  assign t[166] = ~(x[7] & t[187]);
  assign t[167] = t[392] ? t[124] : t[166];
  assign t[168] = ~(t[175] | t[127]);
  assign t[169] = t[392] ? t[188] : t[166];
  assign t[16] = ~(t[392] & t[393]);
  assign t[170] = ~(t[430]);
  assign t[171] = ~(t[422] | t[423]);
  assign t[172] = ~(t[81] | t[189]);
  assign t[173] = t[395] & t[190];
  assign t[174] = ~(t[191]);
  assign t[175] = ~(t[81] | t[192]);
  assign t[176] = ~(t[193] & t[191]);
  assign t[177] = ~(t[81] | t[194]);
  assign t[178] = ~(t[79] & t[195]);
  assign t[179] = ~(t[173] & t[196]);
  assign t[17] = ~(t[394] & t[395]);
  assign t[180] = ~(t[431]);
  assign t[181] = ~(t[427] | t[428]);
  assign t[182] = t[184] | t[131];
  assign t[183] = ~(t[197] & t[85]);
  assign t[184] = ~(t[191] & t[198]);
  assign t[185] = ~(t[393]);
  assign t[186] = ~(t[159] & t[395]);
  assign t[187] = ~(t[393] | t[395]);
  assign t[188] = ~(t[395] & t[163]);
  assign t[189] = t[392] ? t[166] : t[188];
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[79] | t[392]);
  assign t[191] = ~(t[199] | t[129]);
  assign t[192] = t[392] ? t[123] : t[124];
  assign t[193] = ~(t[126] | t[146]);
  assign t[194] = t[392] ? t[122] : t[186];
  assign t[195] = ~(t[166] & t[188]);
  assign t[196] = t[161] | t[159];
  assign t[197] = ~(t[200] | t[175]);
  assign t[198] = ~(t[162] & t[201]);
  assign t[199] = ~(t[79] | t[202]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[203]);
  assign t[201] = t[81] & t[392];
  assign t[202] = t[392] ? t[121] : t[122];
  assign t[203] = ~(t[190] & t[204]);
  assign t[204] = ~(t[188] & t[123]);
  assign t[205] = t[1] ? t[206] : t[432];
  assign t[206] = x[6] ? t[208] : t[207];
  assign t[207] = x[7] ? t[210] : t[209];
  assign t[208] = t[211] ^ x[117];
  assign t[209] = t[212] ^ t[213];
  assign t[20] = t[30] ? x[9] : x[10];
  assign t[210] = ~(t[214] ^ t[215]);
  assign t[211] = x[118] ^ x[119];
  assign t[212] = t[30] ? x[118] : x[119];
  assign t[213] = ~(t[216] ^ t[217]);
  assign t[214] = x[7] ? t[219] : t[218];
  assign t[215] = ~(t[220] ^ t[221]);
  assign t[216] = x[7] ? t[223] : t[222];
  assign t[217] = ~(t[224] ^ t[225]);
  assign t[218] = ~(t[226] & t[227]);
  assign t[219] = t[228] ^ t[218];
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = x[7] ? t[230] : t[229];
  assign t[221] = x[7] ? t[232] : t[231];
  assign t[222] = ~(t[233] & t[234]);
  assign t[223] = t[235] ^ t[236];
  assign t[224] = x[7] ? t[238] : t[237];
  assign t[225] = x[7] ? t[240] : t[239];
  assign t[226] = ~(t[398] & t[54]);
  assign t[227] = ~(t[407] & t[241]);
  assign t[228] = t[88] ? x[121] : x[120];
  assign t[229] = ~(t[242] & t[243]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = t[244] ^ t[237];
  assign t[231] = ~(t[245] & t[246]);
  assign t[232] = t[247] ^ t[248];
  assign t[233] = ~(t[402] & t[66]);
  assign t[234] = ~(t[413] & t[249]);
  assign t[235] = t[88] ? x[123] : x[122];
  assign t[236] = ~(t[250] & t[251]);
  assign t[237] = ~(t[252] & t[253]);
  assign t[238] = t[254] ^ t[239];
  assign t[239] = ~(t[255] & t[256]);
  assign t[23] = ~(t[22] ^ t[35]);
  assign t[240] = t[257] ^ t[258];
  assign t[241] = ~(t[399] & t[53]);
  assign t[242] = ~(t[411] & t[99]);
  assign t[243] = ~(t[424] & t[259]);
  assign t[244] = t[141] ? x[125] : x[124];
  assign t[245] = ~(t[408] & t[92]);
  assign t[246] = ~(t[421] & t[260]);
  assign t[247] = t[88] ? x[127] : x[126];
  assign t[248] = ~(t[261] & t[262]);
  assign t[249] = ~(t[403] & t[65]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = ~(t[414] & t[106]);
  assign t[251] = ~(t[425] & t[263]);
  assign t[252] = ~(t[419] & t[117]);
  assign t[253] = ~(t[429] & t[264]);
  assign t[254] = t[141] ? x[129] : x[128];
  assign t[255] = ~(t[416] & t[110]);
  assign t[256] = ~(t[426] & t[265]);
  assign t[257] = t[30] ? x[131] : x[130];
  assign t[258] = ~(t[266] & t[267]);
  assign t[259] = ~(t[412] & t[98]);
  assign t[25] = x[7] ? t[39] : t[38];
  assign t[260] = ~(t[409] & t[91]);
  assign t[261] = ~(t[422] & t[135]);
  assign t[262] = ~(t[430] & t[268]);
  assign t[263] = ~(t[415] & t[105]);
  assign t[264] = ~(t[420] & t[116]);
  assign t[265] = ~(t[417] & t[109]);
  assign t[266] = ~(t[427] & t[151]);
  assign t[267] = ~(t[431] & t[269]);
  assign t[268] = ~(t[423] & t[134]);
  assign t[269] = ~(t[428] & t[150]);
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[1] ? t[271] : t[433];
  assign t[271] = x[6] ? t[273] : t[272];
  assign t[272] = x[7] ? t[275] : t[274];
  assign t[273] = t[276] ^ x[133];
  assign t[274] = t[277] ^ t[278];
  assign t[275] = ~(t[279] ^ t[280]);
  assign t[276] = x[134] ^ x[135];
  assign t[277] = t[141] ? x[134] : x[135];
  assign t[278] = ~(t[281] ^ t[282]);
  assign t[279] = x[7] ? t[284] : t[283];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = ~(t[285] ^ t[286]);
  assign t[281] = x[7] ? t[288] : t[287];
  assign t[282] = ~(t[289] ^ t[290]);
  assign t[283] = ~(t[291] & t[292]);
  assign t[284] = t[293] ^ t[283];
  assign t[285] = x[7] ? t[295] : t[294];
  assign t[286] = x[7] ? t[297] : t[296];
  assign t[287] = ~(t[298] & t[299]);
  assign t[288] = t[300] ^ t[301];
  assign t[289] = x[7] ? t[303] : t[302];
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = x[7] ? t[305] : t[304];
  assign t[291] = ~(t[54] & t[86]);
  assign t[292] = ~(t[306] & t[396]);
  assign t[293] = t[88] ? x[137] : x[136];
  assign t[294] = ~(t[307] & t[308]);
  assign t[295] = t[309] ^ t[304];
  assign t[296] = ~(t[310] & t[311]);
  assign t[297] = t[312] ^ t[313];
  assign t[298] = ~(t[66] & t[103]);
  assign t[299] = ~(t[314] & t[397]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[30] ? x[139] : x[138];
  assign t[301] = ~(t[315] & t[316]);
  assign t[302] = ~(t[317] & t[318]);
  assign t[303] = t[319] ^ t[320];
  assign t[304] = ~(t[321] & t[322]);
  assign t[305] = t[323] ^ t[302];
  assign t[306] = ~(t[324] & t[53]);
  assign t[307] = ~(t[99] & t[139]);
  assign t[308] = ~(t[325] & t[401]);
  assign t[309] = t[141] ? x[141] : x[140];
  assign t[30] = ~(t[48]);
  assign t[310] = ~(t[92] & t[132]);
  assign t[311] = ~(t[326] & t[400]);
  assign t[312] = t[88] ? x[143] : x[142];
  assign t[313] = ~(t[327] & t[328]);
  assign t[314] = ~(t[329] & t[65]);
  assign t[315] = ~(t[106] & t[144]);
  assign t[316] = ~(t[330] & t[404]);
  assign t[317] = ~(t[110] & t[148]);
  assign t[318] = ~(t[331] & t[405]);
  assign t[319] = t[30] ? x[145] : x[144];
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = ~(t[332] & t[333]);
  assign t[321] = ~(t[117] & t[155]);
  assign t[322] = ~(t[334] & t[406]);
  assign t[323] = t[394] ? x[147] : x[146];
  assign t[324] = ~(t[407] & t[399]);
  assign t[325] = ~(t[335] & t[98]);
  assign t[326] = ~(t[336] & t[91]);
  assign t[327] = ~(t[135] & t[170]);
  assign t[328] = ~(t[337] & t[410]);
  assign t[329] = ~(t[413] & t[403]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = ~(t[338] & t[105]);
  assign t[331] = ~(t[339] & t[109]);
  assign t[332] = ~(t[151] & t[180]);
  assign t[333] = ~(t[340] & t[418]);
  assign t[334] = ~(t[341] & t[116]);
  assign t[335] = ~(t[424] & t[412]);
  assign t[336] = ~(t[421] & t[409]);
  assign t[337] = ~(t[342] & t[134]);
  assign t[338] = ~(t[425] & t[415]);
  assign t[339] = ~(t[426] & t[417]);
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = ~(t[343] & t[150]);
  assign t[341] = ~(t[429] & t[420]);
  assign t[342] = ~(t[430] & t[423]);
  assign t[343] = ~(t[431] & t[428]);
  assign t[344] = t[1] ? t[345] : t[434];
  assign t[345] = x[6] ? t[347] : t[346];
  assign t[346] = x[7] ? t[349] : t[348];
  assign t[347] = t[350] ^ x[149];
  assign t[348] = t[351] ^ t[352];
  assign t[349] = ~(t[353] ^ t[354]);
  assign t[34] = ~(t[396] | t[55]);
  assign t[350] = x[150] ^ x[151];
  assign t[351] = t[88] ? x[150] : x[151];
  assign t[352] = ~(t[355] ^ t[356]);
  assign t[353] = x[7] ? t[358] : t[357];
  assign t[354] = ~(t[359] ^ t[360]);
  assign t[355] = x[7] ? t[362] : t[361];
  assign t[356] = ~(t[363] ^ t[364]);
  assign t[357] = ~(t[291] & t[365]);
  assign t[358] = t[366] ^ t[357];
  assign t[359] = x[7] ? t[368] : t[367];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = x[7] ? t[370] : t[369];
  assign t[361] = ~(t[298] & t[371]);
  assign t[362] = t[372] ^ t[373];
  assign t[363] = x[7] ? t[375] : t[374];
  assign t[364] = x[7] ? t[377] : t[376];
  assign t[365] = t[33] | t[396];
  assign t[366] = t[88] ? x[153] : x[152];
  assign t[367] = ~(t[307] & t[378]);
  assign t[368] = t[379] ^ t[376];
  assign t[369] = ~(t[310] & t[380]);
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[381] ^ t[382];
  assign t[371] = t[40] | t[397];
  assign t[372] = t[30] ? x[155] : x[154];
  assign t[373] = ~(t[315] & t[383]);
  assign t[374] = ~(t[317] & t[384]);
  assign t[375] = t[385] ^ t[386];
  assign t[376] = ~(t[321] & t[387]);
  assign t[377] = t[388] ^ t[374];
  assign t[378] = t[62] | t[401];
  assign t[379] = t[141] ? x[157] : x[156];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[380] = t[58] | t[400];
  assign t[381] = t[88] ? x[159] : x[158];
  assign t[382] = ~(t[327] & t[389]);
  assign t[383] = t[68] | t[404];
  assign t[384] = t[72] | t[405];
  assign t[385] = t[30] ? x[161] : x[160];
  assign t[386] = ~(t[332] & t[390]);
  assign t[387] = t[76] | t[406];
  assign t[388] = t[30] ? x[163] : x[162];
  assign t[389] = t[94] | t[410];
  assign t[38] = ~(t[62] | t[63]);
  assign t[390] = t[112] | t[418];
  assign t[391] = (t[435]);
  assign t[392] = (t[436]);
  assign t[393] = (t[437]);
  assign t[394] = (t[438]);
  assign t[395] = (t[439]);
  assign t[396] = (t[440]);
  assign t[397] = (t[441]);
  assign t[398] = (t[442]);
  assign t[399] = (t[443]);
  assign t[39] = ~(t[46] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (t[444]);
  assign t[401] = (t[445]);
  assign t[402] = (t[446]);
  assign t[403] = (t[447]);
  assign t[404] = (t[448]);
  assign t[405] = (t[449]);
  assign t[406] = (t[450]);
  assign t[407] = (t[451]);
  assign t[408] = (t[452]);
  assign t[409] = (t[453]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (t[454]);
  assign t[411] = (t[455]);
  assign t[412] = (t[456]);
  assign t[413] = (t[457]);
  assign t[414] = (t[458]);
  assign t[415] = (t[459]);
  assign t[416] = (t[460]);
  assign t[417] = (t[461]);
  assign t[418] = (t[462]);
  assign t[419] = (t[463]);
  assign t[41] = ~(t[397] | t[67]);
  assign t[420] = (t[464]);
  assign t[421] = (t[465]);
  assign t[422] = (t[466]);
  assign t[423] = (t[467]);
  assign t[424] = (t[468]);
  assign t[425] = (t[469]);
  assign t[426] = (t[470]);
  assign t[427] = (t[471]);
  assign t[428] = (t[472]);
  assign t[429] = (t[473]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (t[474]);
  assign t[431] = (t[475]);
  assign t[432] = (t[476]);
  assign t[433] = (t[477]);
  assign t[434] = (t[478]);
  assign t[435] = t[479] ^ x[5];
  assign t[436] = t[480] ^ x[13];
  assign t[437] = t[481] ^ x[16];
  assign t[438] = t[482] ^ x[19];
  assign t[439] = t[483] ^ x[22];
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = t[484] ^ x[28];
  assign t[441] = t[485] ^ x[34];
  assign t[442] = t[486] ^ x[35];
  assign t[443] = t[487] ^ x[36];
  assign t[444] = t[488] ^ x[44];
  assign t[445] = t[489] ^ x[50];
  assign t[446] = t[490] ^ x[51];
  assign t[447] = t[491] ^ x[52];
  assign t[448] = t[492] ^ x[58];
  assign t[449] = t[493] ^ x[66];
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = t[494] ^ x[72];
  assign t[451] = t[495] ^ x[73];
  assign t[452] = t[496] ^ x[74];
  assign t[453] = t[497] ^ x[75];
  assign t[454] = t[498] ^ x[81];
  assign t[455] = t[499] ^ x[84];
  assign t[456] = t[500] ^ x[85];
  assign t[457] = t[501] ^ x[88];
  assign t[458] = t[502] ^ x[89];
  assign t[459] = t[503] ^ x[90];
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[460] = t[504] ^ x[91];
  assign t[461] = t[505] ^ x[92];
  assign t[462] = t[506] ^ x[98];
  assign t[463] = t[507] ^ x[101];
  assign t[464] = t[508] ^ x[102];
  assign t[465] = t[509] ^ x[105];
  assign t[466] = t[510] ^ x[106];
  assign t[467] = t[511] ^ x[107];
  assign t[468] = t[512] ^ x[108];
  assign t[469] = t[513] ^ x[109];
  assign t[46] = ~(t[76] | t[77]);
  assign t[470] = t[514] ^ x[110];
  assign t[471] = t[515] ^ x[111];
  assign t[472] = t[516] ^ x[112];
  assign t[473] = t[517] ^ x[113];
  assign t[474] = t[518] ^ x[114];
  assign t[475] = t[519] ^ x[115];
  assign t[476] = t[520] ^ x[116];
  assign t[477] = t[521] ^ x[132];
  assign t[478] = t[522] ^ x[148];
  assign t[479] = (~t[523] & t[524]);
  assign t[47] = ~(t[44] ^ t[78]);
  assign t[480] = (~t[525] & t[526]);
  assign t[481] = (~t[527] & t[528]);
  assign t[482] = (~t[529] & t[530]);
  assign t[483] = (~t[531] & t[532]);
  assign t[484] = (~t[533] & t[534]);
  assign t[485] = (~t[535] & t[536]);
  assign t[486] = (~t[533] & t[537]);
  assign t[487] = (~t[533] & t[538]);
  assign t[488] = (~t[539] & t[540]);
  assign t[489] = (~t[541] & t[542]);
  assign t[48] = ~(t[394]);
  assign t[490] = (~t[535] & t[543]);
  assign t[491] = (~t[535] & t[544]);
  assign t[492] = (~t[545] & t[546]);
  assign t[493] = (~t[547] & t[548]);
  assign t[494] = (~t[549] & t[550]);
  assign t[495] = (~t[533] & t[551]);
  assign t[496] = (~t[539] & t[552]);
  assign t[497] = (~t[539] & t[553]);
  assign t[498] = (~t[554] & t[555]);
  assign t[499] = (~t[541] & t[556]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[541] & t[557]);
  assign t[501] = (~t[535] & t[558]);
  assign t[502] = (~t[545] & t[559]);
  assign t[503] = (~t[545] & t[560]);
  assign t[504] = (~t[547] & t[561]);
  assign t[505] = (~t[547] & t[562]);
  assign t[506] = (~t[563] & t[564]);
  assign t[507] = (~t[549] & t[565]);
  assign t[508] = (~t[549] & t[566]);
  assign t[509] = (~t[539] & t[567]);
  assign t[50] = ~(t[81] | t[82]);
  assign t[510] = (~t[554] & t[568]);
  assign t[511] = (~t[554] & t[569]);
  assign t[512] = (~t[541] & t[570]);
  assign t[513] = (~t[545] & t[571]);
  assign t[514] = (~t[547] & t[572]);
  assign t[515] = (~t[563] & t[573]);
  assign t[516] = (~t[563] & t[574]);
  assign t[517] = (~t[549] & t[575]);
  assign t[518] = (~t[554] & t[576]);
  assign t[519] = (~t[563] & t[577]);
  assign t[51] = ~(t[81] | t[83]);
  assign t[520] = (~t[523] & t[578]);
  assign t[521] = (~t[523] & t[579]);
  assign t[522] = (~t[523] & t[580]);
  assign t[523] = t[581] ^ x[4];
  assign t[524] = t[582] ^ x[5];
  assign t[525] = t[583] ^ x[12];
  assign t[526] = t[584] ^ x[13];
  assign t[527] = t[585] ^ x[15];
  assign t[528] = t[586] ^ x[16];
  assign t[529] = t[587] ^ x[18];
  assign t[52] = ~(t[84] & t[85]);
  assign t[530] = t[588] ^ x[19];
  assign t[531] = t[589] ^ x[21];
  assign t[532] = t[590] ^ x[22];
  assign t[533] = t[591] ^ x[27];
  assign t[534] = t[592] ^ x[28];
  assign t[535] = t[593] ^ x[33];
  assign t[536] = t[594] ^ x[34];
  assign t[537] = t[595] ^ x[35];
  assign t[538] = t[596] ^ x[36];
  assign t[539] = t[597] ^ x[43];
  assign t[53] = ~(t[398]);
  assign t[540] = t[598] ^ x[44];
  assign t[541] = t[599] ^ x[49];
  assign t[542] = t[600] ^ x[50];
  assign t[543] = t[601] ^ x[51];
  assign t[544] = t[602] ^ x[52];
  assign t[545] = t[603] ^ x[57];
  assign t[546] = t[604] ^ x[58];
  assign t[547] = t[605] ^ x[65];
  assign t[548] = t[606] ^ x[66];
  assign t[549] = t[607] ^ x[71];
  assign t[54] = ~(t[399]);
  assign t[550] = t[608] ^ x[72];
  assign t[551] = t[609] ^ x[73];
  assign t[552] = t[610] ^ x[74];
  assign t[553] = t[611] ^ x[75];
  assign t[554] = t[612] ^ x[80];
  assign t[555] = t[613] ^ x[81];
  assign t[556] = t[614] ^ x[84];
  assign t[557] = t[615] ^ x[85];
  assign t[558] = t[616] ^ x[88];
  assign t[559] = t[617] ^ x[89];
  assign t[55] = ~(t[86] | t[87]);
  assign t[560] = t[618] ^ x[90];
  assign t[561] = t[619] ^ x[91];
  assign t[562] = t[620] ^ x[92];
  assign t[563] = t[621] ^ x[97];
  assign t[564] = t[622] ^ x[98];
  assign t[565] = t[623] ^ x[101];
  assign t[566] = t[624] ^ x[102];
  assign t[567] = t[625] ^ x[105];
  assign t[568] = t[626] ^ x[106];
  assign t[569] = t[627] ^ x[107];
  assign t[56] = t[88] ? x[38] : x[37];
  assign t[570] = t[628] ^ x[108];
  assign t[571] = t[629] ^ x[109];
  assign t[572] = t[630] ^ x[110];
  assign t[573] = t[631] ^ x[111];
  assign t[574] = t[632] ^ x[112];
  assign t[575] = t[633] ^ x[113];
  assign t[576] = t[634] ^ x[114];
  assign t[577] = t[635] ^ x[115];
  assign t[578] = t[636] ^ x[116];
  assign t[579] = t[637] ^ x[132];
  assign t[57] = ~(t[89] & t[90]);
  assign t[580] = t[638] ^ x[148];
  assign t[581] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[582] = (x[0]);
  assign t[583] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[584] = (x[11]);
  assign t[585] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[586] = (x[14]);
  assign t[587] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[588] = (x[17]);
  assign t[589] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = ~(t[91] | t[92]);
  assign t[590] = (x[20]);
  assign t[591] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[592] = (x[24]);
  assign t[593] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[594] = (x[30]);
  assign t[595] = (x[25]);
  assign t[596] = (x[26]);
  assign t[597] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[598] = (x[40]);
  assign t[599] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[59] = ~(t[400] | t[93]);
  assign t[5] = t[9] ^ x[8];
  assign t[600] = (x[46]);
  assign t[601] = (x[31]);
  assign t[602] = (x[32]);
  assign t[603] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[604] = (x[54]);
  assign t[605] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[606] = (x[62]);
  assign t[607] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[608] = (x[68]);
  assign t[609] = (x[23]);
  assign t[60] = ~(t[94] | t[95]);
  assign t[610] = (x[41]);
  assign t[611] = (x[42]);
  assign t[612] = (x[76] & ~x[77] & ~x[78] & ~x[79]) | (~x[76] & x[77] & ~x[78] & ~x[79]) | (~x[76] & ~x[77] & x[78] & ~x[79]) | (~x[76] & ~x[77] & ~x[78] & x[79]) | (x[76] & x[77] & x[78] & ~x[79]) | (x[76] & x[77] & ~x[78] & x[79]) | (x[76] & ~x[77] & x[78] & x[79]) | (~x[76] & x[77] & x[78] & x[79]);
  assign t[613] = (x[77]);
  assign t[614] = (x[47]);
  assign t[615] = (x[48]);
  assign t[616] = (x[29]);
  assign t[617] = (x[55]);
  assign t[618] = (x[56]);
  assign t[619] = (x[63]);
  assign t[61] = ~(t[96] ^ t[97]);
  assign t[620] = (x[64]);
  assign t[621] = (x[93] & ~x[94] & ~x[95] & ~x[96]) | (~x[93] & x[94] & ~x[95] & ~x[96]) | (~x[93] & ~x[94] & x[95] & ~x[96]) | (~x[93] & ~x[94] & ~x[95] & x[96]) | (x[93] & x[94] & x[95] & ~x[96]) | (x[93] & x[94] & ~x[95] & x[96]) | (x[93] & ~x[94] & x[95] & x[96]) | (~x[93] & x[94] & x[95] & x[96]);
  assign t[622] = (x[94]);
  assign t[623] = (x[69]);
  assign t[624] = (x[70]);
  assign t[625] = (x[39]);
  assign t[626] = (x[78]);
  assign t[627] = (x[79]);
  assign t[628] = (x[45]);
  assign t[629] = (x[53]);
  assign t[62] = ~(t[98] | t[99]);
  assign t[630] = (x[61]);
  assign t[631] = (x[95]);
  assign t[632] = (x[96]);
  assign t[633] = (x[67]);
  assign t[634] = (x[76]);
  assign t[635] = (x[93]);
  assign t[636] = (x[1]);
  assign t[637] = (x[2]);
  assign t[638] = (x[3]);
  assign t[63] = ~(t[401] | t[100]);
  assign t[64] = ~(t[101] ^ t[102]);
  assign t[65] = ~(t[402]);
  assign t[66] = ~(t[403]);
  assign t[67] = ~(t[103] | t[104]);
  assign t[68] = ~(t[105] | t[106]);
  assign t[69] = ~(t[404] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[30] ? x[60] : x[59];
  assign t[71] = ~(t[108] & t[84]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[405] | t[111]);
  assign t[74] = ~(t[112] | t[113]);
  assign t[75] = ~(t[114] ^ t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[406] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[394]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[392] ? t[122] : t[121];
  assign t[81] = ~(t[79]);
  assign t[82] = t[392] ? t[124] : t[123];
  assign t[83] = t[392] ? t[125] : t[121];
  assign t[84] = ~(t[126] | t[127]);
  assign t[85] = t[79] | t[128];
  assign t[86] = ~(t[407]);
  assign t[87] = ~(t[398] | t[399]);
  assign t[88] = ~(t[48]);
  assign t[89] = ~(t[49] | t[129]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[130] | t[131]);
  assign t[91] = ~(t[408]);
  assign t[92] = ~(t[409]);
  assign t[93] = ~(t[132] | t[133]);
  assign t[94] = ~(t[134] | t[135]);
  assign t[95] = ~(t[410] | t[136]);
  assign t[96] = t[88] ? x[83] : x[82];
  assign t[97] = ~(t[137] & t[138]);
  assign t[98] = ~(t[411]);
  assign t[99] = ~(t[412]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[205] & ~t[270] & ~t[344]) | (~t[0] & t[205] & ~t[270] & ~t[344]) | (~t[0] & ~t[205] & t[270] & ~t[344]) | (~t[0] & ~t[205] & ~t[270] & t[344]) | (t[0] & t[205] & t[270] & ~t[344]) | (t[0] & t[205] & ~t[270] & t[344]) | (t[0] & ~t[205] & t[270] & t[344]) | (~t[0] & t[205] & t[270] & t[344]);
endmodule

module R2ind136(x, y);
 input [115:0] x;
 output y;

 wire [335:0] t;
  assign t[0] = t[1] ? t[2] : t[103];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = ~(t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = t[185] ^ x[5];
  assign t[145] = t[186] ^ x[13];
  assign t[146] = t[187] ^ x[16];
  assign t[147] = t[188] ^ x[19];
  assign t[148] = t[189] ^ x[22];
  assign t[149] = t[190] ^ x[28];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[36];
  assign t[151] = t[192] ^ x[39];
  assign t[152] = t[193] ^ x[40];
  assign t[153] = t[194] ^ x[46];
  assign t[154] = t[195] ^ x[54];
  assign t[155] = t[196] ^ x[57];
  assign t[156] = t[197] ^ x[58];
  assign t[157] = t[198] ^ x[64];
  assign t[158] = t[199] ^ x[70];
  assign t[159] = t[200] ^ x[78];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[81];
  assign t[161] = t[202] ^ x[82];
  assign t[162] = t[203] ^ x[83];
  assign t[163] = t[204] ^ x[84];
  assign t[164] = t[205] ^ x[85];
  assign t[165] = t[206] ^ x[91];
  assign t[166] = t[207] ^ x[92];
  assign t[167] = t[208] ^ x[93];
  assign t[168] = t[209] ^ x[94];
  assign t[169] = t[210] ^ x[95];
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = t[211] ^ x[96];
  assign t[171] = t[212] ^ x[102];
  assign t[172] = t[213] ^ x[103];
  assign t[173] = t[214] ^ x[104];
  assign t[174] = t[215] ^ x[105];
  assign t[175] = t[216] ^ x[106];
  assign t[176] = t[217] ^ x[107];
  assign t[177] = t[218] ^ x[108];
  assign t[178] = t[219] ^ x[109];
  assign t[179] = t[220] ^ x[110];
  assign t[17] = ~(t[106] & t[107]);
  assign t[180] = t[221] ^ x[111];
  assign t[181] = t[222] ^ x[112];
  assign t[182] = t[223] ^ x[113];
  assign t[183] = t[224] ^ x[114];
  assign t[184] = t[225] ^ x[115];
  assign t[185] = (~t[226] & t[227]);
  assign t[186] = (~t[228] & t[229]);
  assign t[187] = (~t[230] & t[231]);
  assign t[188] = (~t[232] & t[233]);
  assign t[189] = (~t[234] & t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = (~t[236] & t[237]);
  assign t[191] = (~t[238] & t[239]);
  assign t[192] = (~t[236] & t[240]);
  assign t[193] = (~t[236] & t[241]);
  assign t[194] = (~t[242] & t[243]);
  assign t[195] = (~t[244] & t[245]);
  assign t[196] = (~t[238] & t[246]);
  assign t[197] = (~t[238] & t[247]);
  assign t[198] = (~t[248] & t[249]);
  assign t[199] = (~t[250] & t[251]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[252] & t[253]);
  assign t[201] = (~t[236] & t[254]);
  assign t[202] = (~t[242] & t[255]);
  assign t[203] = (~t[242] & t[256]);
  assign t[204] = (~t[244] & t[257]);
  assign t[205] = (~t[244] & t[258]);
  assign t[206] = (~t[259] & t[260]);
  assign t[207] = (~t[238] & t[261]);
  assign t[208] = (~t[248] & t[262]);
  assign t[209] = (~t[248] & t[263]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[250] & t[264]);
  assign t[211] = (~t[250] & t[265]);
  assign t[212] = (~t[266] & t[267]);
  assign t[213] = (~t[252] & t[268]);
  assign t[214] = (~t[252] & t[269]);
  assign t[215] = (~t[242] & t[270]);
  assign t[216] = (~t[244] & t[271]);
  assign t[217] = (~t[259] & t[272]);
  assign t[218] = (~t[259] & t[273]);
  assign t[219] = (~t[248] & t[274]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[250] & t[275]);
  assign t[221] = (~t[266] & t[276]);
  assign t[222] = (~t[266] & t[277]);
  assign t[223] = (~t[252] & t[278]);
  assign t[224] = (~t[259] & t[279]);
  assign t[225] = (~t[266] & t[280]);
  assign t[226] = t[281] ^ x[4];
  assign t[227] = t[282] ^ x[5];
  assign t[228] = t[283] ^ x[12];
  assign t[229] = t[284] ^ x[13];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[285] ^ x[15];
  assign t[231] = t[286] ^ x[16];
  assign t[232] = t[287] ^ x[18];
  assign t[233] = t[288] ^ x[19];
  assign t[234] = t[289] ^ x[21];
  assign t[235] = t[290] ^ x[22];
  assign t[236] = t[291] ^ x[27];
  assign t[237] = t[292] ^ x[28];
  assign t[238] = t[293] ^ x[35];
  assign t[239] = t[294] ^ x[36];
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = t[295] ^ x[39];
  assign t[241] = t[296] ^ x[40];
  assign t[242] = t[297] ^ x[45];
  assign t[243] = t[298] ^ x[46];
  assign t[244] = t[299] ^ x[53];
  assign t[245] = t[300] ^ x[54];
  assign t[246] = t[301] ^ x[57];
  assign t[247] = t[302] ^ x[58];
  assign t[248] = t[303] ^ x[63];
  assign t[249] = t[304] ^ x[64];
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = t[305] ^ x[69];
  assign t[251] = t[306] ^ x[70];
  assign t[252] = t[307] ^ x[77];
  assign t[253] = t[308] ^ x[78];
  assign t[254] = t[309] ^ x[81];
  assign t[255] = t[310] ^ x[82];
  assign t[256] = t[311] ^ x[83];
  assign t[257] = t[312] ^ x[84];
  assign t[258] = t[313] ^ x[85];
  assign t[259] = t[314] ^ x[90];
  assign t[25] = ~(t[106]);
  assign t[260] = t[315] ^ x[91];
  assign t[261] = t[316] ^ x[92];
  assign t[262] = t[317] ^ x[93];
  assign t[263] = t[318] ^ x[94];
  assign t[264] = t[319] ^ x[95];
  assign t[265] = t[320] ^ x[96];
  assign t[266] = t[321] ^ x[101];
  assign t[267] = t[322] ^ x[102];
  assign t[268] = t[323] ^ x[103];
  assign t[269] = t[324] ^ x[104];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[325] ^ x[105];
  assign t[271] = t[326] ^ x[106];
  assign t[272] = t[327] ^ x[107];
  assign t[273] = t[328] ^ x[108];
  assign t[274] = t[329] ^ x[109];
  assign t[275] = t[330] ^ x[110];
  assign t[276] = t[331] ^ x[111];
  assign t[277] = t[332] ^ x[112];
  assign t[278] = t[333] ^ x[113];
  assign t[279] = t[334] ^ x[114];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[335] ^ x[115];
  assign t[281] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[282] = (x[3]);
  assign t[283] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[284] = (x[11]);
  assign t[285] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[286] = (x[14]);
  assign t[287] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[288] = (x[17]);
  assign t[289] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[290] = (x[20]);
  assign t[291] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[292] = (x[24]);
  assign t[293] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[294] = (x[32]);
  assign t[295] = (x[26]);
  assign t[296] = (x[23]);
  assign t[297] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[298] = (x[42]);
  assign t[299] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[50]);
  assign t[301] = (x[34]);
  assign t[302] = (x[31]);
  assign t[303] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[304] = (x[60]);
  assign t[305] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[306] = (x[66]);
  assign t[307] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[308] = (x[74]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[44]);
  assign t[311] = (x[41]);
  assign t[312] = (x[52]);
  assign t[313] = (x[49]);
  assign t[314] = (x[86] & ~x[87] & ~x[88] & ~x[89]) | (~x[86] & x[87] & ~x[88] & ~x[89]) | (~x[86] & ~x[87] & x[88] & ~x[89]) | (~x[86] & ~x[87] & ~x[88] & x[89]) | (x[86] & x[87] & x[88] & ~x[89]) | (x[86] & x[87] & ~x[88] & x[89]) | (x[86] & ~x[87] & x[88] & x[89]) | (~x[86] & x[87] & x[88] & x[89]);
  assign t[315] = (x[87]);
  assign t[316] = (x[33]);
  assign t[317] = (x[62]);
  assign t[318] = (x[59]);
  assign t[319] = (x[68]);
  assign t[31] = t[47] | t[108];
  assign t[320] = (x[65]);
  assign t[321] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[322] = (x[98]);
  assign t[323] = (x[76]);
  assign t[324] = (x[73]);
  assign t[325] = (x[43]);
  assign t[326] = (x[51]);
  assign t[327] = (x[89]);
  assign t[328] = (x[86]);
  assign t[329] = (x[61]);
  assign t[32] = t[18] ? x[30] : x[29];
  assign t[330] = (x[67]);
  assign t[331] = (x[100]);
  assign t[332] = (x[97]);
  assign t[333] = (x[75]);
  assign t[334] = (x[88]);
  assign t[335] = (x[99]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] ^ t[43];
  assign t[35] = ~(t[51] & t[52]);
  assign t[36] = t[53] ^ t[54];
  assign t[37] = ~(t[55] & t[56]);
  assign t[38] = t[57] | t[109];
  assign t[39] = t[58] ? x[38] : x[37];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[64];
  assign t[43] = ~(t[65] & t[66]);
  assign t[44] = t[67] ^ t[41];
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[111]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = t[71] | t[112];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[72] ? x[48] : x[47];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = t[75] | t[113];
  assign t[53] = t[18] ? x[56] : x[55];
  assign t[54] = ~(t[76] & t[77]);
  assign t[55] = ~(t[114]);
  assign t[56] = ~(t[115]);
  assign t[57] = ~(t[78] | t[55]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[79] & t[80]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[81] | t[116];
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = t[84] | t[117];
  assign t[63] = t[58] ? x[72] : x[71];
  assign t[64] = ~(t[85] & t[86]);
  assign t[65] = ~(t[87] & t[88]);
  assign t[66] = t[89] | t[118];
  assign t[67] = t[58] ? x[80] : x[79];
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[121]);
  assign t[71] = ~(t[90] | t[69]);
  assign t[72] = ~(t[25]);
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[123]);
  assign t[75] = ~(t[91] | t[73]);
  assign t[76] = ~(t[92] & t[93]);
  assign t[77] = t[94] | t[124];
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[95] | t[79]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[129]);
  assign t[84] = ~(t[96] | t[82]);
  assign t[85] = ~(t[97] & t[98]);
  assign t[86] = t[99] | t[130];
  assign t[87] = ~(t[131]);
  assign t[88] = ~(t[132]);
  assign t[89] = ~(t[100] | t[87]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[136]);
  assign t[94] = ~(t[101] | t[92]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[102] | t[97]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [115:0] x;
 output y;

 wire [344:0] t;
  assign t[0] = t[1] ? t[2] : t[112];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[138] & t[137]);
  assign t[102] = ~(t[147]);
  assign t[103] = ~(t[148]);
  assign t[104] = ~(t[149]);
  assign t[105] = ~(t[110] & t[111]);
  assign t[106] = ~(t[141] & t[140]);
  assign t[107] = ~(t[150]);
  assign t[108] = ~(t[145] & t[144]);
  assign t[109] = ~(t[151]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[149] & t[148]);
  assign t[111] = ~(t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = t[194] ^ x[5];
  assign t[154] = t[195] ^ x[13];
  assign t[155] = t[196] ^ x[16];
  assign t[156] = t[197] ^ x[19];
  assign t[157] = t[198] ^ x[22];
  assign t[158] = t[199] ^ x[28];
  assign t[159] = t[200] ^ x[36];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[39];
  assign t[161] = t[202] ^ x[40];
  assign t[162] = t[203] ^ x[46];
  assign t[163] = t[204] ^ x[54];
  assign t[164] = t[205] ^ x[57];
  assign t[165] = t[206] ^ x[58];
  assign t[166] = t[207] ^ x[64];
  assign t[167] = t[208] ^ x[70];
  assign t[168] = t[209] ^ x[78];
  assign t[169] = t[210] ^ x[81];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[82];
  assign t[171] = t[212] ^ x[83];
  assign t[172] = t[213] ^ x[84];
  assign t[173] = t[214] ^ x[85];
  assign t[174] = t[215] ^ x[91];
  assign t[175] = t[216] ^ x[92];
  assign t[176] = t[217] ^ x[93];
  assign t[177] = t[218] ^ x[94];
  assign t[178] = t[219] ^ x[95];
  assign t[179] = t[220] ^ x[96];
  assign t[17] = ~(t[115] & t[116]);
  assign t[180] = t[221] ^ x[102];
  assign t[181] = t[222] ^ x[103];
  assign t[182] = t[223] ^ x[104];
  assign t[183] = t[224] ^ x[105];
  assign t[184] = t[225] ^ x[106];
  assign t[185] = t[226] ^ x[107];
  assign t[186] = t[227] ^ x[108];
  assign t[187] = t[228] ^ x[109];
  assign t[188] = t[229] ^ x[110];
  assign t[189] = t[230] ^ x[111];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[112];
  assign t[191] = t[232] ^ x[113];
  assign t[192] = t[233] ^ x[114];
  assign t[193] = t[234] ^ x[115];
  assign t[194] = (~t[235] & t[236]);
  assign t[195] = (~t[237] & t[238]);
  assign t[196] = (~t[239] & t[240]);
  assign t[197] = (~t[241] & t[242]);
  assign t[198] = (~t[243] & t[244]);
  assign t[199] = (~t[245] & t[246]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[247] & t[248]);
  assign t[201] = (~t[245] & t[249]);
  assign t[202] = (~t[245] & t[250]);
  assign t[203] = (~t[251] & t[252]);
  assign t[204] = (~t[253] & t[254]);
  assign t[205] = (~t[247] & t[255]);
  assign t[206] = (~t[247] & t[256]);
  assign t[207] = (~t[257] & t[258]);
  assign t[208] = (~t[259] & t[260]);
  assign t[209] = (~t[261] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[245] & t[263]);
  assign t[211] = (~t[251] & t[264]);
  assign t[212] = (~t[251] & t[265]);
  assign t[213] = (~t[253] & t[266]);
  assign t[214] = (~t[253] & t[267]);
  assign t[215] = (~t[268] & t[269]);
  assign t[216] = (~t[247] & t[270]);
  assign t[217] = (~t[257] & t[271]);
  assign t[218] = (~t[257] & t[272]);
  assign t[219] = (~t[259] & t[273]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[259] & t[274]);
  assign t[221] = (~t[275] & t[276]);
  assign t[222] = (~t[261] & t[277]);
  assign t[223] = (~t[261] & t[278]);
  assign t[224] = (~t[251] & t[279]);
  assign t[225] = (~t[253] & t[280]);
  assign t[226] = (~t[268] & t[281]);
  assign t[227] = (~t[268] & t[282]);
  assign t[228] = (~t[257] & t[283]);
  assign t[229] = (~t[259] & t[284]);
  assign t[22] = t[32] ^ t[21];
  assign t[230] = (~t[275] & t[285]);
  assign t[231] = (~t[275] & t[286]);
  assign t[232] = (~t[261] & t[287]);
  assign t[233] = (~t[268] & t[288]);
  assign t[234] = (~t[275] & t[289]);
  assign t[235] = t[290] ^ x[4];
  assign t[236] = t[291] ^ x[5];
  assign t[237] = t[292] ^ x[12];
  assign t[238] = t[293] ^ x[13];
  assign t[239] = t[294] ^ x[15];
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = t[295] ^ x[16];
  assign t[241] = t[296] ^ x[18];
  assign t[242] = t[297] ^ x[19];
  assign t[243] = t[298] ^ x[21];
  assign t[244] = t[299] ^ x[22];
  assign t[245] = t[300] ^ x[27];
  assign t[246] = t[301] ^ x[28];
  assign t[247] = t[302] ^ x[35];
  assign t[248] = t[303] ^ x[36];
  assign t[249] = t[304] ^ x[39];
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = t[305] ^ x[40];
  assign t[251] = t[306] ^ x[45];
  assign t[252] = t[307] ^ x[46];
  assign t[253] = t[308] ^ x[53];
  assign t[254] = t[309] ^ x[54];
  assign t[255] = t[310] ^ x[57];
  assign t[256] = t[311] ^ x[58];
  assign t[257] = t[312] ^ x[63];
  assign t[258] = t[313] ^ x[64];
  assign t[259] = t[314] ^ x[69];
  assign t[25] = ~(t[115]);
  assign t[260] = t[315] ^ x[70];
  assign t[261] = t[316] ^ x[77];
  assign t[262] = t[317] ^ x[78];
  assign t[263] = t[318] ^ x[81];
  assign t[264] = t[319] ^ x[82];
  assign t[265] = t[320] ^ x[83];
  assign t[266] = t[321] ^ x[84];
  assign t[267] = t[322] ^ x[85];
  assign t[268] = t[323] ^ x[90];
  assign t[269] = t[324] ^ x[91];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[325] ^ x[92];
  assign t[271] = t[326] ^ x[93];
  assign t[272] = t[327] ^ x[94];
  assign t[273] = t[328] ^ x[95];
  assign t[274] = t[329] ^ x[96];
  assign t[275] = t[330] ^ x[101];
  assign t[276] = t[331] ^ x[102];
  assign t[277] = t[332] ^ x[103];
  assign t[278] = t[333] ^ x[104];
  assign t[279] = t[334] ^ x[105];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[335] ^ x[106];
  assign t[281] = t[336] ^ x[107];
  assign t[282] = t[337] ^ x[108];
  assign t[283] = t[338] ^ x[109];
  assign t[284] = t[339] ^ x[110];
  assign t[285] = t[340] ^ x[111];
  assign t[286] = t[341] ^ x[112];
  assign t[287] = t[342] ^ x[113];
  assign t[288] = t[343] ^ x[114];
  assign t[289] = t[344] ^ x[115];
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[290] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[291] = (x[2]);
  assign t[292] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[293] = (x[11]);
  assign t[294] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[295] = (x[14]);
  assign t[296] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[297] = (x[17]);
  assign t[298] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[299] = (x[20]);
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[301] = (x[24]);
  assign t[302] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[303] = (x[32]);
  assign t[304] = (x[26]);
  assign t[305] = (x[23]);
  assign t[306] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[307] = (x[42]);
  assign t[308] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[309] = (x[50]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[34]);
  assign t[311] = (x[31]);
  assign t[312] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[313] = (x[60]);
  assign t[314] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[315] = (x[66]);
  assign t[316] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[317] = (x[74]);
  assign t[318] = (x[25]);
  assign t[319] = (x[44]);
  assign t[31] = ~(t[47] & t[117]);
  assign t[320] = (x[41]);
  assign t[321] = (x[52]);
  assign t[322] = (x[49]);
  assign t[323] = (x[86] & ~x[87] & ~x[88] & ~x[89]) | (~x[86] & x[87] & ~x[88] & ~x[89]) | (~x[86] & ~x[87] & x[88] & ~x[89]) | (~x[86] & ~x[87] & ~x[88] & x[89]) | (x[86] & x[87] & x[88] & ~x[89]) | (x[86] & x[87] & ~x[88] & x[89]) | (x[86] & ~x[87] & x[88] & x[89]) | (~x[86] & x[87] & x[88] & x[89]);
  assign t[324] = (x[87]);
  assign t[325] = (x[33]);
  assign t[326] = (x[62]);
  assign t[327] = (x[59]);
  assign t[328] = (x[68]);
  assign t[329] = (x[65]);
  assign t[32] = t[48] ? x[30] : x[29];
  assign t[330] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[331] = (x[98]);
  assign t[332] = (x[76]);
  assign t[333] = (x[73]);
  assign t[334] = (x[43]);
  assign t[335] = (x[51]);
  assign t[336] = (x[89]);
  assign t[337] = (x[86]);
  assign t[338] = (x[61]);
  assign t[339] = (x[67]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[100]);
  assign t[341] = (x[97]);
  assign t[342] = (x[75]);
  assign t[343] = (x[88]);
  assign t[344] = (x[99]);
  assign t[34] = t[51] ^ t[43];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[55];
  assign t[37] = ~(t[56] & t[57]);
  assign t[38] = ~(t[58] & t[118]);
  assign t[39] = t[59] ? x[38] : x[37];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = t[64] ^ t[65];
  assign t[43] = ~(t[66] & t[67]);
  assign t[44] = t[68] ^ t[41];
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[120]);
  assign t[47] = ~(t[69] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[121]);
  assign t[51] = t[18] ? x[48] : x[47];
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = ~(t[76] & t[122]);
  assign t[54] = t[48] ? x[56] : x[55];
  assign t[55] = ~(t[77] & t[78]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[124]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[25]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = ~(t[83] & t[125]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = ~(t[86] & t[126]);
  assign t[64] = t[59] ? x[72] : x[71];
  assign t[65] = ~(t[87] & t[88]);
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = ~(t[91] & t[127]);
  assign t[68] = t[115] ? x[80] : x[79];
  assign t[69] = ~(t[120] & t[119]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[130]);
  assign t[73] = ~(t[92] & t[93]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[132]);
  assign t[76] = ~(t[94] & t[95]);
  assign t[77] = ~(t[96] & t[97]);
  assign t[78] = ~(t[98] & t[133]);
  assign t[79] = ~(t[124] & t[123]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[99] & t[100]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[138]);
  assign t[86] = ~(t[101] & t[102]);
  assign t[87] = ~(t[103] & t[104]);
  assign t[88] = ~(t[105] & t[139]);
  assign t[89] = ~(t[140]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[141]);
  assign t[91] = ~(t[106] & t[107]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[132] & t[131]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[144]);
  assign t[97] = ~(t[145]);
  assign t[98] = ~(t[108] & t[109]);
  assign t[99] = ~(t[136] & t[135]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [106:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[5];
  assign t[127] = t[159] ^ x[13];
  assign t[128] = t[160] ^ x[16];
  assign t[129] = t[161] ^ x[19];
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = t[162] ^ x[22];
  assign t[131] = t[163] ^ x[28];
  assign t[132] = t[164] ^ x[29];
  assign t[133] = t[165] ^ x[37];
  assign t[134] = t[166] ^ x[38];
  assign t[135] = t[167] ^ x[41];
  assign t[136] = t[168] ^ x[47];
  assign t[137] = t[169] ^ x[48];
  assign t[138] = t[170] ^ x[56];
  assign t[139] = t[171] ^ x[57];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[60];
  assign t[141] = t[173] ^ x[66];
  assign t[142] = t[174] ^ x[67];
  assign t[143] = t[175] ^ x[73];
  assign t[144] = t[176] ^ x[74];
  assign t[145] = t[177] ^ x[82];
  assign t[146] = t[178] ^ x[83];
  assign t[147] = t[179] ^ x[86];
  assign t[148] = t[180] ^ x[87];
  assign t[149] = t[181] ^ x[93];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[94];
  assign t[151] = t[183] ^ x[95];
  assign t[152] = t[184] ^ x[96];
  assign t[153] = t[185] ^ x[97];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[104];
  assign t[156] = t[188] ^ x[105];
  assign t[157] = t[189] ^ x[106];
  assign t[158] = (~t[190] & t[191]);
  assign t[159] = (~t[192] & t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (~t[194] & t[195]);
  assign t[161] = (~t[196] & t[197]);
  assign t[162] = (~t[198] & t[199]);
  assign t[163] = (~t[200] & t[201]);
  assign t[164] = (~t[200] & t[202]);
  assign t[165] = (~t[203] & t[204]);
  assign t[166] = (~t[203] & t[205]);
  assign t[167] = (~t[200] & t[206]);
  assign t[168] = (~t[207] & t[208]);
  assign t[169] = (~t[207] & t[209]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (~t[210] & t[211]);
  assign t[171] = (~t[210] & t[212]);
  assign t[172] = (~t[203] & t[213]);
  assign t[173] = (~t[214] & t[215]);
  assign t[174] = (~t[214] & t[216]);
  assign t[175] = (~t[217] & t[218]);
  assign t[176] = (~t[217] & t[219]);
  assign t[177] = (~t[220] & t[221]);
  assign t[178] = (~t[220] & t[222]);
  assign t[179] = (~t[207] & t[223]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (~t[210] & t[224]);
  assign t[181] = (~t[225] & t[226]);
  assign t[182] = (~t[225] & t[227]);
  assign t[183] = (~t[214] & t[228]);
  assign t[184] = (~t[217] & t[229]);
  assign t[185] = (~t[220] & t[230]);
  assign t[186] = (~t[231] & t[232]);
  assign t[187] = (~t[231] & t[233]);
  assign t[188] = (~t[225] & t[234]);
  assign t[189] = (~t[231] & t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[236] ^ x[4];
  assign t[191] = t[237] ^ x[5];
  assign t[192] = t[238] ^ x[12];
  assign t[193] = t[239] ^ x[13];
  assign t[194] = t[240] ^ x[15];
  assign t[195] = t[241] ^ x[16];
  assign t[196] = t[242] ^ x[18];
  assign t[197] = t[243] ^ x[19];
  assign t[198] = t[244] ^ x[21];
  assign t[199] = t[245] ^ x[22];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[246] ^ x[27];
  assign t[201] = t[247] ^ x[28];
  assign t[202] = t[248] ^ x[29];
  assign t[203] = t[249] ^ x[36];
  assign t[204] = t[250] ^ x[37];
  assign t[205] = t[251] ^ x[38];
  assign t[206] = t[252] ^ x[41];
  assign t[207] = t[253] ^ x[46];
  assign t[208] = t[254] ^ x[47];
  assign t[209] = t[255] ^ x[48];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[256] ^ x[55];
  assign t[211] = t[257] ^ x[56];
  assign t[212] = t[258] ^ x[57];
  assign t[213] = t[259] ^ x[60];
  assign t[214] = t[260] ^ x[65];
  assign t[215] = t[261] ^ x[66];
  assign t[216] = t[262] ^ x[67];
  assign t[217] = t[263] ^ x[72];
  assign t[218] = t[264] ^ x[73];
  assign t[219] = t[265] ^ x[74];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[266] ^ x[81];
  assign t[221] = t[267] ^ x[82];
  assign t[222] = t[268] ^ x[83];
  assign t[223] = t[269] ^ x[86];
  assign t[224] = t[270] ^ x[87];
  assign t[225] = t[271] ^ x[92];
  assign t[226] = t[272] ^ x[93];
  assign t[227] = t[273] ^ x[94];
  assign t[228] = t[274] ^ x[95];
  assign t[229] = t[275] ^ x[96];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[276] ^ x[97];
  assign t[231] = t[277] ^ x[102];
  assign t[232] = t[278] ^ x[103];
  assign t[233] = t[279] ^ x[104];
  assign t[234] = t[280] ^ x[105];
  assign t[235] = t[281] ^ x[106];
  assign t[236] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[237] = (x[1]);
  assign t[238] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[239] = (x[11]);
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[241] = (x[14]);
  assign t[242] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[243] = (x[17]);
  assign t[244] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[245] = (x[20]);
  assign t[246] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[247] = (x[25]);
  assign t[248] = (x[23]);
  assign t[249] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = (x[34]);
  assign t[251] = (x[32]);
  assign t[252] = (x[26]);
  assign t[253] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[254] = (x[44]);
  assign t[255] = (x[42]);
  assign t[256] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[257] = (x[53]);
  assign t[258] = (x[51]);
  assign t[259] = (x[35]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[261] = (x[63]);
  assign t[262] = (x[61]);
  assign t[263] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[264] = (x[70]);
  assign t[265] = (x[68]);
  assign t[266] = (x[77] & ~x[78] & ~x[79] & ~x[80]) | (~x[77] & x[78] & ~x[79] & ~x[80]) | (~x[77] & ~x[78] & x[79] & ~x[80]) | (~x[77] & ~x[78] & ~x[79] & x[80]) | (x[77] & x[78] & x[79] & ~x[80]) | (x[77] & x[78] & ~x[79] & x[80]) | (x[77] & ~x[78] & x[79] & x[80]) | (~x[77] & x[78] & x[79] & x[80]);
  assign t[267] = (x[79]);
  assign t[268] = (x[77]);
  assign t[269] = (x[45]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[54]);
  assign t[271] = (x[88] & ~x[89] & ~x[90] & ~x[91]) | (~x[88] & x[89] & ~x[90] & ~x[91]) | (~x[88] & ~x[89] & x[90] & ~x[91]) | (~x[88] & ~x[89] & ~x[90] & x[91]) | (x[88] & x[89] & x[90] & ~x[91]) | (x[88] & x[89] & ~x[90] & x[91]) | (x[88] & ~x[89] & x[90] & x[91]) | (~x[88] & x[89] & x[90] & x[91]);
  assign t[272] = (x[90]);
  assign t[273] = (x[88]);
  assign t[274] = (x[64]);
  assign t[275] = (x[71]);
  assign t[276] = (x[80]);
  assign t[277] = (x[98] & ~x[99] & ~x[100] & ~x[101]) | (~x[98] & x[99] & ~x[100] & ~x[101]) | (~x[98] & ~x[99] & x[100] & ~x[101]) | (~x[98] & ~x[99] & ~x[100] & x[101]) | (x[98] & x[99] & x[100] & ~x[101]) | (x[98] & x[99] & ~x[100] & x[101]) | (x[98] & ~x[99] & x[100] & x[101]) | (~x[98] & x[99] & x[100] & x[101]);
  assign t[278] = (x[100]);
  assign t[279] = (x[98]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[91]);
  assign t[281] = (x[101]);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[47] ? x[31] : x[30];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] ^ t[41];
  assign t[35] = ~(t[51] & t[52]);
  assign t[36] = t[53] ^ t[54];
  assign t[37] = ~(t[101] & t[55]);
  assign t[38] = ~(t[102] & t[56]);
  assign t[39] = t[47] ? x[40] : x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = t[61] ^ t[43];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[65];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[66]);
  assign t[47] = ~(t[25]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = ~(t[105] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[69] ? x[50] : x[49];
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = t[47] ? x[59] : x[58];
  assign t[54] = ~(t[72] & t[73]);
  assign t[55] = ~(t[108]);
  assign t[56] = ~(t[108] & t[74]);
  assign t[57] = ~(t[109] & t[75]);
  assign t[58] = ~(t[110] & t[76]);
  assign t[59] = ~(t[111] & t[77]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[112] & t[78]);
  assign t[61] = t[69] ? x[76] : x[75];
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = ~(t[114] & t[80]);
  assign t[64] = t[18] ? x[85] : x[84];
  assign t[65] = ~(t[81] & t[82]);
  assign t[66] = ~(t[99]);
  assign t[67] = ~(t[115]);
  assign t[68] = ~(t[115] & t[83]);
  assign t[69] = ~(t[25]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[116]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[117] & t[85]);
  assign t[73] = ~(t[118] & t[86]);
  assign t[74] = ~(t[101]);
  assign t[75] = ~(t[119]);
  assign t[76] = ~(t[119] & t[87]);
  assign t[77] = ~(t[120]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[106]);
  assign t[85] = ~(t[124]);
  assign t[86] = ~(t[124] & t[92]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125]);
  assign t[91] = ~(t[125] & t[93]);
  assign t[92] = ~(t[117]);
  assign t[93] = ~(t[122]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [115:0] x;
 output y;

 wire [437:0] t;
  assign t[0] = t[1] ? t[2] : t[205];
  assign t[100] = ~(t[139] | t[140]);
  assign t[101] = t[141] ? x[87] : x[86];
  assign t[102] = ~(t[142] & t[143]);
  assign t[103] = ~(t[227]);
  assign t[104] = ~(t[216] | t[217]);
  assign t[105] = ~(t[228]);
  assign t[106] = ~(t[229]);
  assign t[107] = ~(t[144] | t[145]);
  assign t[108] = ~(t[146] | t[147]);
  assign t[109] = ~(t[230]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[231]);
  assign t[111] = ~(t[148] | t[149]);
  assign t[112] = ~(t[150] | t[151]);
  assign t[113] = ~(t[232] | t[152]);
  assign t[114] = t[30] ? x[100] : x[99];
  assign t[115] = ~(t[153] & t[154]);
  assign t[116] = ~(t[233]);
  assign t[117] = ~(t[234]);
  assign t[118] = ~(t[155] | t[156]);
  assign t[119] = t[30] ? x[104] : x[103];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[157] & t[158]);
  assign t[121] = ~(t[159] & t[160]);
  assign t[122] = ~(t[161] & t[160]);
  assign t[123] = ~(x[7] & t[162]);
  assign t[124] = ~(t[163] & t[160]);
  assign t[125] = ~(t[161] & t[209]);
  assign t[126] = ~(t[81] | t[164]);
  assign t[127] = ~(t[81] | t[165]);
  assign t[128] = t[206] ? t[166] : t[124];
  assign t[129] = ~(t[79] | t[167]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[168]);
  assign t[131] = ~(t[81] | t[169]);
  assign t[132] = ~(t[235]);
  assign t[133] = ~(t[222] | t[223]);
  assign t[134] = ~(t[236]);
  assign t[135] = ~(t[237]);
  assign t[136] = ~(t[170] | t[171]);
  assign t[137] = ~(t[172] | t[127]);
  assign t[138] = ~(t[173] | t[174]);
  assign t[139] = ~(t[238]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[225] | t[226]);
  assign t[141] = ~(t[48]);
  assign t[142] = ~(t[175] | t[176]);
  assign t[143] = ~(t[177]);
  assign t[144] = ~(t[239]);
  assign t[145] = ~(t[228] | t[229]);
  assign t[146] = ~(t[31] & t[178]);
  assign t[147] = ~(t[179] & t[85]);
  assign t[148] = ~(t[240]);
  assign t[149] = ~(t[230] | t[231]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[241]);
  assign t[151] = ~(t[242]);
  assign t[152] = ~(t[180] | t[181]);
  assign t[153] = ~(t[126] | t[172]);
  assign t[154] = ~(t[182] | t[183]);
  assign t[155] = ~(t[243]);
  assign t[156] = ~(t[233] | t[234]);
  assign t[157] = ~(t[177] | t[51]);
  assign t[158] = ~(t[49] | t[184]);
  assign t[159] = x[7] & t[207];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[209]);
  assign t[161] = ~(x[7] | t[207]);
  assign t[162] = ~(t[207] | t[160]);
  assign t[163] = ~(x[7] | t[185]);
  assign t[164] = t[206] ? t[186] : t[122];
  assign t[165] = t[206] ? t[121] : t[125];
  assign t[166] = ~(x[7] & t[187]);
  assign t[167] = t[206] ? t[124] : t[166];
  assign t[168] = ~(t[175] | t[127]);
  assign t[169] = t[206] ? t[188] : t[166];
  assign t[16] = ~(t[206] & t[207]);
  assign t[170] = ~(t[244]);
  assign t[171] = ~(t[236] | t[237]);
  assign t[172] = ~(t[81] | t[189]);
  assign t[173] = t[209] & t[190];
  assign t[174] = ~(t[191]);
  assign t[175] = ~(t[81] | t[192]);
  assign t[176] = ~(t[193] & t[191]);
  assign t[177] = ~(t[81] | t[194]);
  assign t[178] = ~(t[79] & t[195]);
  assign t[179] = ~(t[173] & t[196]);
  assign t[17] = ~(t[208] & t[209]);
  assign t[180] = ~(t[245]);
  assign t[181] = ~(t[241] | t[242]);
  assign t[182] = t[184] | t[131];
  assign t[183] = ~(t[197] & t[85]);
  assign t[184] = ~(t[191] & t[198]);
  assign t[185] = ~(t[207]);
  assign t[186] = ~(t[159] & t[209]);
  assign t[187] = ~(t[207] | t[209]);
  assign t[188] = ~(t[209] & t[163]);
  assign t[189] = t[206] ? t[166] : t[188];
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[79] | t[206]);
  assign t[191] = ~(t[199] | t[129]);
  assign t[192] = t[206] ? t[123] : t[124];
  assign t[193] = ~(t[126] | t[146]);
  assign t[194] = t[206] ? t[122] : t[186];
  assign t[195] = ~(t[166] & t[188]);
  assign t[196] = t[161] | t[159];
  assign t[197] = ~(t[200] | t[175]);
  assign t[198] = ~(t[162] & t[201]);
  assign t[199] = ~(t[79] | t[202]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[203]);
  assign t[201] = t[81] & t[206];
  assign t[202] = t[206] ? t[121] : t[122];
  assign t[203] = ~(t[190] & t[204]);
  assign t[204] = ~(t[188] & t[123]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[9] : x[10];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[22] ^ t[35]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = (t[283]);
  assign t[243] = (t[284]);
  assign t[244] = (t[285]);
  assign t[245] = (t[286]);
  assign t[246] = t[287] ^ x[5];
  assign t[247] = t[288] ^ x[13];
  assign t[248] = t[289] ^ x[16];
  assign t[249] = t[290] ^ x[19];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[22];
  assign t[251] = t[292] ^ x[28];
  assign t[252] = t[293] ^ x[34];
  assign t[253] = t[294] ^ x[35];
  assign t[254] = t[295] ^ x[36];
  assign t[255] = t[296] ^ x[44];
  assign t[256] = t[297] ^ x[50];
  assign t[257] = t[298] ^ x[51];
  assign t[258] = t[299] ^ x[52];
  assign t[259] = t[300] ^ x[58];
  assign t[25] = x[7] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[66];
  assign t[261] = t[302] ^ x[72];
  assign t[262] = t[303] ^ x[73];
  assign t[263] = t[304] ^ x[74];
  assign t[264] = t[305] ^ x[75];
  assign t[265] = t[306] ^ x[81];
  assign t[266] = t[307] ^ x[84];
  assign t[267] = t[308] ^ x[85];
  assign t[268] = t[309] ^ x[88];
  assign t[269] = t[310] ^ x[89];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[90];
  assign t[271] = t[312] ^ x[91];
  assign t[272] = t[313] ^ x[92];
  assign t[273] = t[314] ^ x[98];
  assign t[274] = t[315] ^ x[101];
  assign t[275] = t[316] ^ x[102];
  assign t[276] = t[317] ^ x[105];
  assign t[277] = t[318] ^ x[106];
  assign t[278] = t[319] ^ x[107];
  assign t[279] = t[320] ^ x[108];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[321] ^ x[109];
  assign t[281] = t[322] ^ x[110];
  assign t[282] = t[323] ^ x[111];
  assign t[283] = t[324] ^ x[112];
  assign t[284] = t[325] ^ x[113];
  assign t[285] = t[326] ^ x[114];
  assign t[286] = t[327] ^ x[115];
  assign t[287] = (~t[328] & t[329]);
  assign t[288] = (~t[330] & t[331]);
  assign t[289] = (~t[332] & t[333]);
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = (~t[334] & t[335]);
  assign t[291] = (~t[336] & t[337]);
  assign t[292] = (~t[338] & t[339]);
  assign t[293] = (~t[340] & t[341]);
  assign t[294] = (~t[338] & t[342]);
  assign t[295] = (~t[338] & t[343]);
  assign t[296] = (~t[344] & t[345]);
  assign t[297] = (~t[346] & t[347]);
  assign t[298] = (~t[340] & t[348]);
  assign t[299] = (~t[340] & t[349]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[350] & t[351]);
  assign t[301] = (~t[352] & t[353]);
  assign t[302] = (~t[354] & t[355]);
  assign t[303] = (~t[338] & t[356]);
  assign t[304] = (~t[344] & t[357]);
  assign t[305] = (~t[344] & t[358]);
  assign t[306] = (~t[359] & t[360]);
  assign t[307] = (~t[346] & t[361]);
  assign t[308] = (~t[346] & t[362]);
  assign t[309] = (~t[340] & t[363]);
  assign t[30] = ~(t[48]);
  assign t[310] = (~t[350] & t[364]);
  assign t[311] = (~t[350] & t[365]);
  assign t[312] = (~t[352] & t[366]);
  assign t[313] = (~t[352] & t[367]);
  assign t[314] = (~t[368] & t[369]);
  assign t[315] = (~t[354] & t[370]);
  assign t[316] = (~t[354] & t[371]);
  assign t[317] = (~t[344] & t[372]);
  assign t[318] = (~t[359] & t[373]);
  assign t[319] = (~t[359] & t[374]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (~t[346] & t[375]);
  assign t[321] = (~t[350] & t[376]);
  assign t[322] = (~t[352] & t[377]);
  assign t[323] = (~t[368] & t[378]);
  assign t[324] = (~t[368] & t[379]);
  assign t[325] = (~t[354] & t[380]);
  assign t[326] = (~t[359] & t[381]);
  assign t[327] = (~t[368] & t[382]);
  assign t[328] = t[383] ^ x[4];
  assign t[329] = t[384] ^ x[5];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[385] ^ x[12];
  assign t[331] = t[386] ^ x[13];
  assign t[332] = t[387] ^ x[15];
  assign t[333] = t[388] ^ x[16];
  assign t[334] = t[389] ^ x[18];
  assign t[335] = t[390] ^ x[19];
  assign t[336] = t[391] ^ x[21];
  assign t[337] = t[392] ^ x[22];
  assign t[338] = t[393] ^ x[27];
  assign t[339] = t[394] ^ x[28];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[395] ^ x[33];
  assign t[341] = t[396] ^ x[34];
  assign t[342] = t[397] ^ x[35];
  assign t[343] = t[398] ^ x[36];
  assign t[344] = t[399] ^ x[43];
  assign t[345] = t[400] ^ x[44];
  assign t[346] = t[401] ^ x[49];
  assign t[347] = t[402] ^ x[50];
  assign t[348] = t[403] ^ x[51];
  assign t[349] = t[404] ^ x[52];
  assign t[34] = ~(t[210] | t[55]);
  assign t[350] = t[405] ^ x[57];
  assign t[351] = t[406] ^ x[58];
  assign t[352] = t[407] ^ x[65];
  assign t[353] = t[408] ^ x[66];
  assign t[354] = t[409] ^ x[71];
  assign t[355] = t[410] ^ x[72];
  assign t[356] = t[411] ^ x[73];
  assign t[357] = t[412] ^ x[74];
  assign t[358] = t[413] ^ x[75];
  assign t[359] = t[414] ^ x[80];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[415] ^ x[81];
  assign t[361] = t[416] ^ x[84];
  assign t[362] = t[417] ^ x[85];
  assign t[363] = t[418] ^ x[88];
  assign t[364] = t[419] ^ x[89];
  assign t[365] = t[420] ^ x[90];
  assign t[366] = t[421] ^ x[91];
  assign t[367] = t[422] ^ x[92];
  assign t[368] = t[423] ^ x[97];
  assign t[369] = t[424] ^ x[98];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[425] ^ x[101];
  assign t[371] = t[426] ^ x[102];
  assign t[372] = t[427] ^ x[105];
  assign t[373] = t[428] ^ x[106];
  assign t[374] = t[429] ^ x[107];
  assign t[375] = t[430] ^ x[108];
  assign t[376] = t[431] ^ x[109];
  assign t[377] = t[432] ^ x[110];
  assign t[378] = t[433] ^ x[111];
  assign t[379] = t[434] ^ x[112];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[380] = t[435] ^ x[113];
  assign t[381] = t[436] ^ x[114];
  assign t[382] = t[437] ^ x[115];
  assign t[383] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[384] = (x[0]);
  assign t[385] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[386] = (x[11]);
  assign t[387] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[388] = (x[14]);
  assign t[389] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = ~(t[62] | t[63]);
  assign t[390] = (x[17]);
  assign t[391] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[392] = (x[20]);
  assign t[393] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[394] = (x[24]);
  assign t[395] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[396] = (x[30]);
  assign t[397] = (x[25]);
  assign t[398] = (x[26]);
  assign t[399] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[39] = ~(t[46] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[40]);
  assign t[401] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[402] = (x[46]);
  assign t[403] = (x[31]);
  assign t[404] = (x[32]);
  assign t[405] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[406] = (x[54]);
  assign t[407] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[408] = (x[62]);
  assign t[409] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[68]);
  assign t[411] = (x[23]);
  assign t[412] = (x[41]);
  assign t[413] = (x[42]);
  assign t[414] = (x[76] & ~x[77] & ~x[78] & ~x[79]) | (~x[76] & x[77] & ~x[78] & ~x[79]) | (~x[76] & ~x[77] & x[78] & ~x[79]) | (~x[76] & ~x[77] & ~x[78] & x[79]) | (x[76] & x[77] & x[78] & ~x[79]) | (x[76] & x[77] & ~x[78] & x[79]) | (x[76] & ~x[77] & x[78] & x[79]) | (~x[76] & x[77] & x[78] & x[79]);
  assign t[415] = (x[77]);
  assign t[416] = (x[47]);
  assign t[417] = (x[48]);
  assign t[418] = (x[29]);
  assign t[419] = (x[55]);
  assign t[41] = ~(t[211] | t[67]);
  assign t[420] = (x[56]);
  assign t[421] = (x[63]);
  assign t[422] = (x[64]);
  assign t[423] = (x[93] & ~x[94] & ~x[95] & ~x[96]) | (~x[93] & x[94] & ~x[95] & ~x[96]) | (~x[93] & ~x[94] & x[95] & ~x[96]) | (~x[93] & ~x[94] & ~x[95] & x[96]) | (x[93] & x[94] & x[95] & ~x[96]) | (x[93] & x[94] & ~x[95] & x[96]) | (x[93] & ~x[94] & x[95] & x[96]) | (~x[93] & x[94] & x[95] & x[96]);
  assign t[424] = (x[94]);
  assign t[425] = (x[69]);
  assign t[426] = (x[70]);
  assign t[427] = (x[39]);
  assign t[428] = (x[78]);
  assign t[429] = (x[79]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[45]);
  assign t[431] = (x[53]);
  assign t[432] = (x[61]);
  assign t[433] = (x[95]);
  assign t[434] = (x[96]);
  assign t[435] = (x[67]);
  assign t[436] = (x[76]);
  assign t[437] = (x[93]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[45] = ~(t[74] ^ t[75]);
  assign t[46] = ~(t[76] | t[77]);
  assign t[47] = ~(t[44] ^ t[78]);
  assign t[48] = ~(t[208]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[81] | t[82]);
  assign t[51] = ~(t[81] | t[83]);
  assign t[52] = ~(t[84] & t[85]);
  assign t[53] = ~(t[212]);
  assign t[54] = ~(t[213]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = t[88] ? x[38] : x[37];
  assign t[57] = ~(t[89] & t[90]);
  assign t[58] = ~(t[91] | t[92]);
  assign t[59] = ~(t[214] | t[93]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[94] | t[95]);
  assign t[61] = ~(t[96] ^ t[97]);
  assign t[62] = ~(t[98] | t[99]);
  assign t[63] = ~(t[215] | t[100]);
  assign t[64] = ~(t[101] ^ t[102]);
  assign t[65] = ~(t[216]);
  assign t[66] = ~(t[217]);
  assign t[67] = ~(t[103] | t[104]);
  assign t[68] = ~(t[105] | t[106]);
  assign t[69] = ~(t[218] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[30] ? x[60] : x[59];
  assign t[71] = ~(t[108] & t[84]);
  assign t[72] = ~(t[109] | t[110]);
  assign t[73] = ~(t[219] | t[111]);
  assign t[74] = ~(t[112] | t[113]);
  assign t[75] = ~(t[114] ^ t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[220] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[208]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[206] ? t[122] : t[121];
  assign t[81] = ~(t[79]);
  assign t[82] = t[206] ? t[124] : t[123];
  assign t[83] = t[206] ? t[125] : t[121];
  assign t[84] = ~(t[126] | t[127]);
  assign t[85] = t[79] | t[128];
  assign t[86] = ~(t[221]);
  assign t[87] = ~(t[212] | t[213]);
  assign t[88] = ~(t[48]);
  assign t[89] = ~(t[49] | t[129]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[130] | t[131]);
  assign t[91] = ~(t[222]);
  assign t[92] = ~(t[223]);
  assign t[93] = ~(t[132] | t[133]);
  assign t[94] = ~(t[134] | t[135]);
  assign t[95] = ~(t[224] | t[136]);
  assign t[96] = t[88] ? x[83] : x[82];
  assign t[97] = ~(t[137] & t[138]);
  assign t[98] = ~(t[225]);
  assign t[99] = ~(t[226]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [112:0] x;
 output y;

 wire [485:0] t;
  assign t[0] = t[1] ? t[2] : t[304];
  assign t[100] = t[63] & t[305];
  assign t[101] = ~(t[327]);
  assign t[102] = ~(t[319] | t[320]);
  assign t[103] = ~(t[328]);
  assign t[104] = ~(t[329]);
  assign t[105] = ~(t[126] | t[127]);
  assign t[106] = ~(t[43] | t[128]);
  assign t[107] = ~(t[42] | t[129]);
  assign t[108] = ~(t[330]);
  assign t[109] = ~(t[322] | t[323]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[331]);
  assign t[111] = ~(t[332]);
  assign t[112] = ~(t[130] | t[131]);
  assign t[113] = ~(t[132] | t[133]);
  assign t[114] = ~(t[117] | t[134]);
  assign t[115] = ~(t[333]);
  assign t[116] = ~(t[325] | t[326]);
  assign t[117] = ~(t[63] | t[135]);
  assign t[118] = ~(t[63] | t[136]);
  assign t[119] = t[44] | t[137];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[138] & t[139]);
  assign t[121] = x[7] & t[306];
  assign t[122] = ~(x[7] | t[306]);
  assign t[123] = ~(t[308]);
  assign t[124] = t[305] ? t[95] : t[94];
  assign t[125] = t[305] ? t[141] : t[140];
  assign t[126] = ~(t[334]);
  assign t[127] = ~(t[328] | t[329]);
  assign t[128] = ~(t[63] | t[142]);
  assign t[129] = ~(t[114] & t[139]);
  assign t[12] = ~(t[18] ^ t[15]);
  assign t[130] = ~(t[335]);
  assign t[131] = ~(t[331] | t[332]);
  assign t[132] = ~(t[106] & t[143]);
  assign t[133] = ~(t[144] & t[139]);
  assign t[134] = ~(t[63] | t[145]);
  assign t[135] = t[305] ? t[93] : t[94];
  assign t[136] = t[305] ? t[140] : t[146];
  assign t[137] = ~(t[63] | t[147]);
  assign t[138] = ~(t[148] | t[149]);
  assign t[139] = t[66] | t[150];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = ~(x[7] & t[151]);
  assign t[141] = ~(t[152] & t[123]);
  assign t[142] = t[305] ? t[141] : t[153];
  assign t[143] = ~(t[66] & t[154]);
  assign t[144] = ~(t[155] & t[156]);
  assign t[145] = t[305] ? t[95] : t[96];
  assign t[146] = ~(t[308] & t[152]);
  assign t[147] = t[305] ? t[146] : t[140];
  assign t[148] = ~(t[157]);
  assign t[149] = ~(t[63] | t[158]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[305] ? t[140] : t[141];
  assign t[151] = ~(t[306] | t[308]);
  assign t[152] = ~(x[7] | t[159]);
  assign t[153] = ~(x[7] & t[99]);
  assign t[154] = ~(t[140] & t[146]);
  assign t[155] = t[308] & t[160];
  assign t[156] = t[122] | t[121];
  assign t[157] = ~(t[160] & t[161]);
  assign t[158] = t[305] ? t[153] : t[141];
  assign t[159] = ~(t[306]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = ~(t[66] | t[305]);
  assign t[161] = ~(t[146] & t[153]);
  assign t[162] = t[1] ? t[163] : t[310];
  assign t[163] = x[6] ? t[165] : t[164];
  assign t[164] = x[7] ? t[167] : t[166];
  assign t[165] = t[168] ^ x[86];
  assign t[166] = t[169] ^ t[170];
  assign t[167] = ~(t[171] ^ t[172]);
  assign t[168] = x[87] ^ x[88];
  assign t[169] = t[173] ? x[87] : x[88];
  assign t[16] = ~(t[305] & t[306]);
  assign t[170] = ~(t[174] ^ t[172]);
  assign t[171] = x[7] ? t[176] : t[175];
  assign t[172] = ~(t[177] ^ t[178]);
  assign t[173] = ~(t[40]);
  assign t[174] = x[7] ? t[180] : t[179];
  assign t[175] = ~(t[181] & t[182]);
  assign t[176] = t[169] ^ t[179];
  assign t[177] = x[7] ? t[184] : t[183];
  assign t[178] = x[7] ? t[186] : t[185];
  assign t[179] = ~(t[187] & t[188]);
  assign t[17] = ~(t[307] & t[308]);
  assign t[180] = t[189] ^ t[190];
  assign t[181] = ~(t[311] & t[46]);
  assign t[182] = ~(t[318] & t[191]);
  assign t[183] = ~(t[192] & t[193]);
  assign t[184] = t[194] ^ t[195];
  assign t[185] = ~(t[196] & t[197]);
  assign t[186] = t[198] ^ t[199];
  assign t[187] = ~(t[315] & t[57]);
  assign t[188] = ~(t[304] & t[200]);
  assign t[189] = t[27] ? x[90] : x[89];
  assign t[18] = x[7] ? t[26] : t[25];
  assign t[190] = ~(t[201] & t[202]);
  assign t[191] = ~(t[312] & t[45]);
  assign t[192] = ~(t[322] & t[80]);
  assign t[193] = ~(t[330] & t[203]);
  assign t[194] = t[204] ? x[92] : x[91];
  assign t[195] = ~(t[205] & t[206]);
  assign t[196] = ~(t[319] & t[73]);
  assign t[197] = ~(t[327] & t[207]);
  assign t[198] = t[27] ? x[94] : x[93];
  assign t[199] = ~(t[208] & t[209]);
  assign t[19] = t[27] ? x[9] : x[10];
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[316] & t[56]);
  assign t[201] = ~(t[325] & t[89]);
  assign t[202] = ~(t[333] & t[210]);
  assign t[203] = ~(t[323] & t[79]);
  assign t[204] = ~(t[40]);
  assign t[205] = ~(t[331] & t[111]);
  assign t[206] = ~(t[335] & t[211]);
  assign t[207] = ~(t[320] & t[72]);
  assign t[208] = ~(t[328] & t[104]);
  assign t[209] = ~(t[334] & t[212]);
  assign t[20] = ~(t[28] & t[29]);
  assign t[210] = ~(t[326] & t[88]);
  assign t[211] = ~(t[332] & t[110]);
  assign t[212] = ~(t[329] & t[103]);
  assign t[213] = t[1] ? t[214] : t[315];
  assign t[214] = x[6] ? t[216] : t[215];
  assign t[215] = x[7] ? t[218] : t[217];
  assign t[216] = t[219] ^ x[95];
  assign t[217] = t[220] ^ t[221];
  assign t[218] = ~(t[222] ^ t[223]);
  assign t[219] = x[96] ^ x[97];
  assign t[21] = ~(t[30] | t[31]);
  assign t[220] = t[307] ? x[96] : x[97];
  assign t[221] = ~(t[224] ^ t[223]);
  assign t[222] = x[7] ? t[226] : t[225];
  assign t[223] = ~(t[227] ^ t[228]);
  assign t[224] = x[7] ? t[230] : t[229];
  assign t[225] = ~(t[231] & t[232]);
  assign t[226] = t[220] ^ t[229];
  assign t[227] = x[7] ? t[234] : t[233];
  assign t[228] = x[7] ? t[236] : t[235];
  assign t[229] = ~(t[237] & t[238]);
  assign t[22] = ~(t[25] ^ t[13]);
  assign t[230] = t[239] ^ t[240];
  assign t[231] = ~(t[46] & t[70]);
  assign t[232] = ~(t[241] & t[309]);
  assign t[233] = ~(t[242] & t[243]);
  assign t[234] = t[244] ^ t[245];
  assign t[235] = ~(t[246] & t[247]);
  assign t[236] = t[248] ^ t[249];
  assign t[237] = ~(t[57] & t[86]);
  assign t[238] = ~(t[250] & t[310]);
  assign t[239] = t[27] ? x[99] : x[98];
  assign t[23] = x[7] ? t[33] : t[32];
  assign t[240] = ~(t[251] & t[252]);
  assign t[241] = ~(t[253] & t[45]);
  assign t[242] = ~(t[80] & t[108]);
  assign t[243] = ~(t[254] & t[314]);
  assign t[244] = t[27] ? x[101] : x[100];
  assign t[245] = ~(t[255] & t[256]);
  assign t[246] = ~(t[73] & t[101]);
  assign t[247] = ~(t[257] & t[313]);
  assign t[248] = t[173] ? x[103] : x[102];
  assign t[249] = ~(t[258] & t[259]);
  assign t[24] = x[7] ? t[35] : t[34];
  assign t[250] = ~(t[260] & t[56]);
  assign t[251] = ~(t[89] & t[115]);
  assign t[252] = ~(t[261] & t[317]);
  assign t[253] = ~(t[318] & t[312]);
  assign t[254] = ~(t[262] & t[79]);
  assign t[255] = ~(t[111] & t[130]);
  assign t[256] = ~(t[263] & t[324]);
  assign t[257] = ~(t[264] & t[72]);
  assign t[258] = ~(t[104] & t[126]);
  assign t[259] = ~(t[265] & t[321]);
  assign t[25] = ~(t[36] | t[37]);
  assign t[260] = ~(t[304] & t[316]);
  assign t[261] = ~(t[266] & t[88]);
  assign t[262] = ~(t[330] & t[323]);
  assign t[263] = ~(t[267] & t[110]);
  assign t[264] = ~(t[327] & t[320]);
  assign t[265] = ~(t[268] & t[103]);
  assign t[266] = ~(t[333] & t[326]);
  assign t[267] = ~(t[335] & t[332]);
  assign t[268] = ~(t[334] & t[329]);
  assign t[269] = t[1] ? t[270] : t[316];
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = x[6] ? t[272] : t[271];
  assign t[271] = x[7] ? t[274] : t[273];
  assign t[272] = t[275] ^ x[104];
  assign t[273] = t[276] ^ t[277];
  assign t[274] = ~(t[278] ^ t[279]);
  assign t[275] = x[105] ^ x[106];
  assign t[276] = t[27] ? x[105] : x[106];
  assign t[277] = ~(t[280] ^ t[279]);
  assign t[278] = x[7] ? t[282] : t[281];
  assign t[279] = ~(t[283] ^ t[284]);
  assign t[27] = ~(t[40]);
  assign t[280] = x[7] ? t[286] : t[285];
  assign t[281] = ~(t[231] & t[287]);
  assign t[282] = t[276] ^ t[285];
  assign t[283] = x[7] ? t[289] : t[288];
  assign t[284] = x[7] ? t[291] : t[290];
  assign t[285] = ~(t[237] & t[292]);
  assign t[286] = t[293] ^ t[294];
  assign t[287] = t[30] | t[309];
  assign t[288] = ~(t[242] & t[295]);
  assign t[289] = t[296] ^ t[297];
  assign t[28] = ~(t[41] | t[42]);
  assign t[290] = ~(t[246] & t[298]);
  assign t[291] = t[299] ^ t[300];
  assign t[292] = t[36] | t[310];
  assign t[293] = t[27] ? x[108] : x[107];
  assign t[294] = ~(t[251] & t[301]);
  assign t[295] = t[52] | t[314];
  assign t[296] = t[27] ? x[110] : x[109];
  assign t[297] = ~(t[255] & t[302]);
  assign t[298] = t[48] | t[313];
  assign t[299] = t[204] ? x[112] : x[111];
  assign t[29] = ~(t[43] | t[44]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = ~(t[258] & t[303]);
  assign t[301] = t[59] | t[317];
  assign t[302] = t[82] | t[324];
  assign t[303] = t[75] | t[321];
  assign t[304] = (t[336]);
  assign t[305] = (t[337]);
  assign t[306] = (t[338]);
  assign t[307] = (t[339]);
  assign t[308] = (t[340]);
  assign t[309] = (t[341]);
  assign t[30] = ~(t[45] | t[46]);
  assign t[310] = (t[342]);
  assign t[311] = (t[343]);
  assign t[312] = (t[344]);
  assign t[313] = (t[345]);
  assign t[314] = (t[346]);
  assign t[315] = (t[347]);
  assign t[316] = (t[348]);
  assign t[317] = (t[349]);
  assign t[318] = (t[350]);
  assign t[319] = (t[351]);
  assign t[31] = ~(t[309] | t[47]);
  assign t[320] = (t[352]);
  assign t[321] = (t[353]);
  assign t[322] = (t[354]);
  assign t[323] = (t[355]);
  assign t[324] = (t[356]);
  assign t[325] = (t[357]);
  assign t[326] = (t[358]);
  assign t[327] = (t[359]);
  assign t[328] = (t[360]);
  assign t[329] = (t[361]);
  assign t[32] = ~(t[48] | t[49]);
  assign t[330] = (t[362]);
  assign t[331] = (t[363]);
  assign t[332] = (t[364]);
  assign t[333] = (t[365]);
  assign t[334] = (t[366]);
  assign t[335] = (t[367]);
  assign t[336] = t[368] ^ x[5];
  assign t[337] = t[369] ^ x[13];
  assign t[338] = t[370] ^ x[16];
  assign t[339] = t[371] ^ x[19];
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[340] = t[372] ^ x[22];
  assign t[341] = t[373] ^ x[28];
  assign t[342] = t[374] ^ x[29];
  assign t[343] = t[375] ^ x[30];
  assign t[344] = t[376] ^ x[31];
  assign t[345] = t[377] ^ x[37];
  assign t[346] = t[378] ^ x[43];
  assign t[347] = t[379] ^ x[44];
  assign t[348] = t[380] ^ x[45];
  assign t[349] = t[381] ^ x[51];
  assign t[34] = ~(t[52] | t[53]);
  assign t[350] = t[382] ^ x[54];
  assign t[351] = t[383] ^ x[55];
  assign t[352] = t[384] ^ x[56];
  assign t[353] = t[385] ^ x[62];
  assign t[354] = t[386] ^ x[65];
  assign t[355] = t[387] ^ x[66];
  assign t[356] = t[388] ^ x[72];
  assign t[357] = t[389] ^ x[75];
  assign t[358] = t[390] ^ x[76];
  assign t[359] = t[391] ^ x[77];
  assign t[35] = ~(t[54] ^ t[55]);
  assign t[360] = t[392] ^ x[78];
  assign t[361] = t[393] ^ x[79];
  assign t[362] = t[394] ^ x[80];
  assign t[363] = t[395] ^ x[81];
  assign t[364] = t[396] ^ x[82];
  assign t[365] = t[397] ^ x[83];
  assign t[366] = t[398] ^ x[84];
  assign t[367] = t[399] ^ x[85];
  assign t[368] = (~t[400] & t[401]);
  assign t[369] = (~t[402] & t[403]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[370] = (~t[404] & t[405]);
  assign t[371] = (~t[406] & t[407]);
  assign t[372] = (~t[408] & t[409]);
  assign t[373] = (~t[410] & t[411]);
  assign t[374] = (~t[400] & t[412]);
  assign t[375] = (~t[410] & t[413]);
  assign t[376] = (~t[410] & t[414]);
  assign t[377] = (~t[415] & t[416]);
  assign t[378] = (~t[417] & t[418]);
  assign t[379] = (~t[400] & t[419]);
  assign t[37] = ~(t[310] | t[58]);
  assign t[380] = (~t[400] & t[420]);
  assign t[381] = (~t[421] & t[422]);
  assign t[382] = (~t[410] & t[423]);
  assign t[383] = (~t[415] & t[424]);
  assign t[384] = (~t[415] & t[425]);
  assign t[385] = (~t[426] & t[427]);
  assign t[386] = (~t[417] & t[428]);
  assign t[387] = (~t[417] & t[429]);
  assign t[388] = (~t[430] & t[431]);
  assign t[389] = (~t[421] & t[432]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[390] = (~t[421] & t[433]);
  assign t[391] = (~t[415] & t[434]);
  assign t[392] = (~t[426] & t[435]);
  assign t[393] = (~t[426] & t[436]);
  assign t[394] = (~t[417] & t[437]);
  assign t[395] = (~t[430] & t[438]);
  assign t[396] = (~t[430] & t[439]);
  assign t[397] = (~t[421] & t[440]);
  assign t[398] = (~t[426] & t[441]);
  assign t[399] = (~t[430] & t[442]);
  assign t[39] = ~(t[61] ^ t[62]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[443] ^ x[4];
  assign t[401] = t[444] ^ x[5];
  assign t[402] = t[445] ^ x[12];
  assign t[403] = t[446] ^ x[13];
  assign t[404] = t[447] ^ x[15];
  assign t[405] = t[448] ^ x[16];
  assign t[406] = t[449] ^ x[18];
  assign t[407] = t[450] ^ x[19];
  assign t[408] = t[451] ^ x[21];
  assign t[409] = t[452] ^ x[22];
  assign t[40] = ~(t[307]);
  assign t[410] = t[453] ^ x[27];
  assign t[411] = t[454] ^ x[28];
  assign t[412] = t[455] ^ x[29];
  assign t[413] = t[456] ^ x[30];
  assign t[414] = t[457] ^ x[31];
  assign t[415] = t[458] ^ x[36];
  assign t[416] = t[459] ^ x[37];
  assign t[417] = t[460] ^ x[42];
  assign t[418] = t[461] ^ x[43];
  assign t[419] = t[462] ^ x[44];
  assign t[41] = ~(t[63] | t[64]);
  assign t[420] = t[463] ^ x[45];
  assign t[421] = t[464] ^ x[50];
  assign t[422] = t[465] ^ x[51];
  assign t[423] = t[466] ^ x[54];
  assign t[424] = t[467] ^ x[55];
  assign t[425] = t[468] ^ x[56];
  assign t[426] = t[469] ^ x[61];
  assign t[427] = t[470] ^ x[62];
  assign t[428] = t[471] ^ x[65];
  assign t[429] = t[472] ^ x[66];
  assign t[42] = ~(t[63] | t[65]);
  assign t[430] = t[473] ^ x[71];
  assign t[431] = t[474] ^ x[72];
  assign t[432] = t[475] ^ x[75];
  assign t[433] = t[476] ^ x[76];
  assign t[434] = t[477] ^ x[77];
  assign t[435] = t[478] ^ x[78];
  assign t[436] = t[479] ^ x[79];
  assign t[437] = t[480] ^ x[80];
  assign t[438] = t[481] ^ x[81];
  assign t[439] = t[482] ^ x[82];
  assign t[43] = ~(t[66] | t[67]);
  assign t[440] = t[483] ^ x[83];
  assign t[441] = t[484] ^ x[84];
  assign t[442] = t[485] ^ x[85];
  assign t[443] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[444] = (x[0]);
  assign t[445] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[446] = (x[11]);
  assign t[447] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[448] = (x[14]);
  assign t[449] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[44] = ~(t[68] & t[69]);
  assign t[450] = (x[17]);
  assign t[451] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[452] = (x[20]);
  assign t[453] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[454] = (x[24]);
  assign t[455] = (x[1]);
  assign t[456] = (x[25]);
  assign t[457] = (x[26]);
  assign t[458] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[459] = (x[33]);
  assign t[45] = ~(t[311]);
  assign t[460] = (x[38] & ~x[39] & ~x[40] & ~x[41]) | (~x[38] & x[39] & ~x[40] & ~x[41]) | (~x[38] & ~x[39] & x[40] & ~x[41]) | (~x[38] & ~x[39] & ~x[40] & x[41]) | (x[38] & x[39] & x[40] & ~x[41]) | (x[38] & x[39] & ~x[40] & x[41]) | (x[38] & ~x[39] & x[40] & x[41]) | (~x[38] & x[39] & x[40] & x[41]);
  assign t[461] = (x[39]);
  assign t[462] = (x[2]);
  assign t[463] = (x[3]);
  assign t[464] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[465] = (x[47]);
  assign t[466] = (x[23]);
  assign t[467] = (x[34]);
  assign t[468] = (x[35]);
  assign t[469] = (x[57] & ~x[58] & ~x[59] & ~x[60]) | (~x[57] & x[58] & ~x[59] & ~x[60]) | (~x[57] & ~x[58] & x[59] & ~x[60]) | (~x[57] & ~x[58] & ~x[59] & x[60]) | (x[57] & x[58] & x[59] & ~x[60]) | (x[57] & x[58] & ~x[59] & x[60]) | (x[57] & ~x[58] & x[59] & x[60]) | (~x[57] & x[58] & x[59] & x[60]);
  assign t[46] = ~(t[312]);
  assign t[470] = (x[58]);
  assign t[471] = (x[40]);
  assign t[472] = (x[41]);
  assign t[473] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[474] = (x[68]);
  assign t[475] = (x[48]);
  assign t[476] = (x[49]);
  assign t[477] = (x[32]);
  assign t[478] = (x[59]);
  assign t[479] = (x[60]);
  assign t[47] = ~(t[70] | t[71]);
  assign t[480] = (x[38]);
  assign t[481] = (x[69]);
  assign t[482] = (x[70]);
  assign t[483] = (x[46]);
  assign t[484] = (x[57]);
  assign t[485] = (x[67]);
  assign t[48] = ~(t[72] | t[73]);
  assign t[49] = ~(t[313] | t[74]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[75] | t[76]);
  assign t[51] = ~(t[77] ^ t[78]);
  assign t[52] = ~(t[79] | t[80]);
  assign t[53] = ~(t[314] | t[81]);
  assign t[54] = ~(t[82] | t[83]);
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = ~(t[315]);
  assign t[57] = ~(t[316]);
  assign t[58] = ~(t[86] | t[87]);
  assign t[59] = ~(t[88] | t[89]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[317] | t[90]);
  assign t[61] = t[27] ? x[53] : x[52];
  assign t[62] = ~(t[91] & t[92]);
  assign t[63] = ~(t[66]);
  assign t[64] = t[305] ? t[94] : t[93];
  assign t[65] = t[305] ? t[96] : t[95];
  assign t[66] = ~(t[307]);
  assign t[67] = t[305] ? t[94] : t[95];
  assign t[68] = ~(t[97] | t[98]);
  assign t[69] = ~(t[99] & t[100]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[318]);
  assign t[71] = ~(t[311] | t[312]);
  assign t[72] = ~(t[319]);
  assign t[73] = ~(t[320]);
  assign t[74] = ~(t[101] | t[102]);
  assign t[75] = ~(t[103] | t[104]);
  assign t[76] = ~(t[321] | t[105]);
  assign t[77] = t[27] ? x[64] : x[63];
  assign t[78] = ~(t[106] & t[107]);
  assign t[79] = ~(t[322]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[323]);
  assign t[81] = ~(t[108] | t[109]);
  assign t[82] = ~(t[110] | t[111]);
  assign t[83] = ~(t[324] | t[112]);
  assign t[84] = t[27] ? x[74] : x[73];
  assign t[85] = ~(t[113] & t[114]);
  assign t[86] = ~(t[304]);
  assign t[87] = ~(t[315] | t[316]);
  assign t[88] = ~(t[325]);
  assign t[89] = ~(t[326]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[115] | t[116]);
  assign t[91] = ~(t[117] | t[118]);
  assign t[92] = ~(t[119] | t[120]);
  assign t[93] = ~(t[121] & t[308]);
  assign t[94] = ~(t[122] & t[123]);
  assign t[95] = ~(t[121] & t[123]);
  assign t[96] = ~(t[122] & t[308]);
  assign t[97] = ~(t[66] | t[124]);
  assign t[98] = ~(t[66] | t[125]);
  assign t[99] = ~(t[306] | t[123]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[162] & ~t[213] & ~t[269]) | (~t[0] & t[162] & ~t[213] & ~t[269]) | (~t[0] & ~t[162] & t[213] & ~t[269]) | (~t[0] & ~t[162] & ~t[213] & t[269]) | (t[0] & t[162] & t[213] & ~t[269]) | (t[0] & t[162] & ~t[213] & t[269]) | (t[0] & ~t[162] & t[213] & t[269]) | (~t[0] & t[162] & t[213] & t[269]);
endmodule

module R2ind141(x, y);
 input [85:0] x;
 output y;

 wire [261:0] t;
  assign t[0] = t[1] ? t[2] : t[80];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = t[144] ^ x[5];
  assign t[113] = t[145] ^ x[13];
  assign t[114] = t[146] ^ x[16];
  assign t[115] = t[147] ^ x[19];
  assign t[116] = t[148] ^ x[22];
  assign t[117] = t[149] ^ x[28];
  assign t[118] = t[150] ^ x[29];
  assign t[119] = t[151] ^ x[32];
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[33];
  assign t[121] = t[153] ^ x[39];
  assign t[122] = t[154] ^ x[47];
  assign t[123] = t[155] ^ x[50];
  assign t[124] = t[156] ^ x[56];
  assign t[125] = t[157] ^ x[57];
  assign t[126] = t[158] ^ x[58];
  assign t[127] = t[159] ^ x[59];
  assign t[128] = t[160] ^ x[65];
  assign t[129] = t[161] ^ x[66];
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = t[162] ^ x[67];
  assign t[131] = t[163] ^ x[73];
  assign t[132] = t[164] ^ x[74];
  assign t[133] = t[165] ^ x[75];
  assign t[134] = t[166] ^ x[76];
  assign t[135] = t[167] ^ x[77];
  assign t[136] = t[168] ^ x[78];
  assign t[137] = t[169] ^ x[79];
  assign t[138] = t[170] ^ x[80];
  assign t[139] = t[171] ^ x[81];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[82];
  assign t[141] = t[173] ^ x[83];
  assign t[142] = t[174] ^ x[84];
  assign t[143] = t[175] ^ x[85];
  assign t[144] = (~t[176] & t[177]);
  assign t[145] = (~t[178] & t[179]);
  assign t[146] = (~t[180] & t[181]);
  assign t[147] = (~t[182] & t[183]);
  assign t[148] = (~t[184] & t[185]);
  assign t[149] = (~t[186] & t[187]);
  assign t[14] = x[7] ? t[21] : t[20];
  assign t[150] = (~t[176] & t[188]);
  assign t[151] = (~t[186] & t[189]);
  assign t[152] = (~t[186] & t[190]);
  assign t[153] = (~t[191] & t[192]);
  assign t[154] = (~t[193] & t[194]);
  assign t[155] = (~t[176] & t[195]);
  assign t[156] = (~t[196] & t[197]);
  assign t[157] = (~t[186] & t[198]);
  assign t[158] = (~t[191] & t[199]);
  assign t[159] = (~t[191] & t[200]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (~t[201] & t[202]);
  assign t[161] = (~t[193] & t[203]);
  assign t[162] = (~t[193] & t[204]);
  assign t[163] = (~t[205] & t[206]);
  assign t[164] = (~t[176] & t[207]);
  assign t[165] = (~t[196] & t[208]);
  assign t[166] = (~t[196] & t[209]);
  assign t[167] = (~t[191] & t[210]);
  assign t[168] = (~t[201] & t[211]);
  assign t[169] = (~t[201] & t[212]);
  assign t[16] = ~(t[81] & t[82]);
  assign t[170] = (~t[193] & t[213]);
  assign t[171] = (~t[205] & t[214]);
  assign t[172] = (~t[205] & t[215]);
  assign t[173] = (~t[196] & t[216]);
  assign t[174] = (~t[201] & t[217]);
  assign t[175] = (~t[205] & t[218]);
  assign t[176] = t[219] ^ x[4];
  assign t[177] = t[220] ^ x[5];
  assign t[178] = t[221] ^ x[12];
  assign t[179] = t[222] ^ x[13];
  assign t[17] = ~(t[83] & t[84]);
  assign t[180] = t[223] ^ x[15];
  assign t[181] = t[224] ^ x[16];
  assign t[182] = t[225] ^ x[18];
  assign t[183] = t[226] ^ x[19];
  assign t[184] = t[227] ^ x[21];
  assign t[185] = t[228] ^ x[22];
  assign t[186] = t[229] ^ x[27];
  assign t[187] = t[230] ^ x[28];
  assign t[188] = t[231] ^ x[29];
  assign t[189] = t[232] ^ x[32];
  assign t[18] = ~(t[24]);
  assign t[190] = t[233] ^ x[33];
  assign t[191] = t[234] ^ x[38];
  assign t[192] = t[235] ^ x[39];
  assign t[193] = t[236] ^ x[46];
  assign t[194] = t[237] ^ x[47];
  assign t[195] = t[238] ^ x[50];
  assign t[196] = t[239] ^ x[55];
  assign t[197] = t[240] ^ x[56];
  assign t[198] = t[241] ^ x[57];
  assign t[199] = t[242] ^ x[58];
  assign t[19] = x[7] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[59];
  assign t[201] = t[244] ^ x[64];
  assign t[202] = t[245] ^ x[65];
  assign t[203] = t[246] ^ x[66];
  assign t[204] = t[247] ^ x[67];
  assign t[205] = t[248] ^ x[72];
  assign t[206] = t[249] ^ x[73];
  assign t[207] = t[250] ^ x[74];
  assign t[208] = t[251] ^ x[75];
  assign t[209] = t[252] ^ x[76];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[253] ^ x[77];
  assign t[211] = t[254] ^ x[78];
  assign t[212] = t[255] ^ x[79];
  assign t[213] = t[256] ^ x[80];
  assign t[214] = t[257] ^ x[81];
  assign t[215] = t[258] ^ x[82];
  assign t[216] = t[259] ^ x[83];
  assign t[217] = t[260] ^ x[84];
  assign t[218] = t[261] ^ x[85];
  assign t[219] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[21] = t[12] ^ t[25];
  assign t[220] = (x[3]);
  assign t[221] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[222] = (x[11]);
  assign t[223] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[224] = (x[14]);
  assign t[225] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[226] = (x[17]);
  assign t[227] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[228] = (x[20]);
  assign t[229] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[22] = x[7] ? t[30] : t[29];
  assign t[230] = (x[24]);
  assign t[231] = (x[1]);
  assign t[232] = (x[26]);
  assign t[233] = (x[23]);
  assign t[234] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[235] = (x[35]);
  assign t[236] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[237] = (x[43]);
  assign t[238] = (x[0]);
  assign t[239] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[23] = x[7] ? t[32] : t[31];
  assign t[240] = (x[52]);
  assign t[241] = (x[25]);
  assign t[242] = (x[37]);
  assign t[243] = (x[34]);
  assign t[244] = (x[60] & ~x[61] & ~x[62] & ~x[63]) | (~x[60] & x[61] & ~x[62] & ~x[63]) | (~x[60] & ~x[61] & x[62] & ~x[63]) | (~x[60] & ~x[61] & ~x[62] & x[63]) | (x[60] & x[61] & x[62] & ~x[63]) | (x[60] & x[61] & ~x[62] & x[63]) | (x[60] & ~x[61] & x[62] & x[63]) | (~x[60] & x[61] & x[62] & x[63]);
  assign t[245] = (x[61]);
  assign t[246] = (x[45]);
  assign t[247] = (x[42]);
  assign t[248] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[249] = (x[69]);
  assign t[24] = ~(t[83]);
  assign t[250] = (x[2]);
  assign t[251] = (x[54]);
  assign t[252] = (x[51]);
  assign t[253] = (x[36]);
  assign t[254] = (x[63]);
  assign t[255] = (x[60]);
  assign t[256] = (x[44]);
  assign t[257] = (x[71]);
  assign t[258] = (x[68]);
  assign t[259] = (x[53]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[62]);
  assign t[261] = (x[70]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[37] & t[38]);
  assign t[28] = t[39] | t[85];
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] | t[86];
  assign t[35] = t[18] ? x[31] : x[30];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[88]);
  assign t[39] = ~(t[53] | t[37]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[89];
  assign t[42] = t[18] ? x[41] : x[40];
  assign t[43] = ~(t[57] & t[58]);
  assign t[44] = ~(t[59] & t[60]);
  assign t[45] = t[61] | t[90];
  assign t[46] = t[62] ? x[49] : x[48];
  assign t[47] = ~(t[63] & t[64]);
  assign t[48] = ~(t[80]);
  assign t[49] = ~(t[91]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[65] | t[48]);
  assign t[51] = ~(t[66] & t[67]);
  assign t[52] = t[68] | t[92];
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[95]);
  assign t[56] = ~(t[69] | t[54]);
  assign t[57] = ~(t[70] & t[71]);
  assign t[58] = t[72] | t[96];
  assign t[59] = ~(t[97]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[98]);
  assign t[61] = ~(t[73] | t[59]);
  assign t[62] = ~(t[24]);
  assign t[63] = ~(t[74] & t[75]);
  assign t[64] = t[76] | t[99];
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[102]);
  assign t[68] = ~(t[77] | t[66]);
  assign t[69] = ~(t[103]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[105]);
  assign t[72] = ~(t[78] | t[70]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[108]);
  assign t[76] = ~(t[79] | t[74]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = ~(t[111]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[112]);
  assign t[81] = (t[113]);
  assign t[82] = (t[114]);
  assign t[83] = (t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [85:0] x;
 output y;

 wire [268:0] t;
  assign t[0] = t[1] ? t[2] : t[87];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = t[151] ^ x[5];
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[13];
  assign t[121] = t[153] ^ x[16];
  assign t[122] = t[154] ^ x[19];
  assign t[123] = t[155] ^ x[22];
  assign t[124] = t[156] ^ x[28];
  assign t[125] = t[157] ^ x[29];
  assign t[126] = t[158] ^ x[32];
  assign t[127] = t[159] ^ x[33];
  assign t[128] = t[160] ^ x[39];
  assign t[129] = t[161] ^ x[47];
  assign t[12] = t[88] ? x[9] : x[10];
  assign t[130] = t[162] ^ x[50];
  assign t[131] = t[163] ^ x[51];
  assign t[132] = t[164] ^ x[57];
  assign t[133] = t[165] ^ x[58];
  assign t[134] = t[166] ^ x[59];
  assign t[135] = t[167] ^ x[60];
  assign t[136] = t[168] ^ x[66];
  assign t[137] = t[169] ^ x[67];
  assign t[138] = t[170] ^ x[68];
  assign t[139] = t[171] ^ x[74];
  assign t[13] = ~(t[18] ^ t[15]);
  assign t[140] = t[172] ^ x[75];
  assign t[141] = t[173] ^ x[76];
  assign t[142] = t[174] ^ x[77];
  assign t[143] = t[175] ^ x[78];
  assign t[144] = t[176] ^ x[79];
  assign t[145] = t[177] ^ x[80];
  assign t[146] = t[178] ^ x[81];
  assign t[147] = t[179] ^ x[82];
  assign t[148] = t[180] ^ x[83];
  assign t[149] = t[181] ^ x[84];
  assign t[14] = x[7] ? t[20] : t[19];
  assign t[150] = t[182] ^ x[85];
  assign t[151] = (~t[183] & t[184]);
  assign t[152] = (~t[185] & t[186]);
  assign t[153] = (~t[187] & t[188]);
  assign t[154] = (~t[189] & t[190]);
  assign t[155] = (~t[191] & t[192]);
  assign t[156] = (~t[193] & t[194]);
  assign t[157] = (~t[183] & t[195]);
  assign t[158] = (~t[193] & t[196]);
  assign t[159] = (~t[193] & t[197]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (~t[198] & t[199]);
  assign t[161] = (~t[200] & t[201]);
  assign t[162] = (~t[183] & t[202]);
  assign t[163] = (~t[183] & t[203]);
  assign t[164] = (~t[204] & t[205]);
  assign t[165] = (~t[193] & t[206]);
  assign t[166] = (~t[198] & t[207]);
  assign t[167] = (~t[198] & t[208]);
  assign t[168] = (~t[209] & t[210]);
  assign t[169] = (~t[200] & t[211]);
  assign t[16] = ~(t[89] & t[90]);
  assign t[170] = (~t[200] & t[212]);
  assign t[171] = (~t[213] & t[214]);
  assign t[172] = (~t[204] & t[215]);
  assign t[173] = (~t[204] & t[216]);
  assign t[174] = (~t[198] & t[217]);
  assign t[175] = (~t[209] & t[218]);
  assign t[176] = (~t[209] & t[219]);
  assign t[177] = (~t[200] & t[220]);
  assign t[178] = (~t[213] & t[221]);
  assign t[179] = (~t[213] & t[222]);
  assign t[17] = ~(t[88] & t[91]);
  assign t[180] = (~t[204] & t[223]);
  assign t[181] = (~t[209] & t[224]);
  assign t[182] = (~t[213] & t[225]);
  assign t[183] = t[226] ^ x[4];
  assign t[184] = t[227] ^ x[5];
  assign t[185] = t[228] ^ x[12];
  assign t[186] = t[229] ^ x[13];
  assign t[187] = t[230] ^ x[15];
  assign t[188] = t[231] ^ x[16];
  assign t[189] = t[232] ^ x[18];
  assign t[18] = x[7] ? t[24] : t[23];
  assign t[190] = t[233] ^ x[19];
  assign t[191] = t[234] ^ x[21];
  assign t[192] = t[235] ^ x[22];
  assign t[193] = t[236] ^ x[27];
  assign t[194] = t[237] ^ x[28];
  assign t[195] = t[238] ^ x[29];
  assign t[196] = t[239] ^ x[32];
  assign t[197] = t[240] ^ x[33];
  assign t[198] = t[241] ^ x[38];
  assign t[199] = t[242] ^ x[39];
  assign t[19] = ~(t[25] & t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[46];
  assign t[201] = t[244] ^ x[47];
  assign t[202] = t[245] ^ x[50];
  assign t[203] = t[246] ^ x[51];
  assign t[204] = t[247] ^ x[56];
  assign t[205] = t[248] ^ x[57];
  assign t[206] = t[249] ^ x[58];
  assign t[207] = t[250] ^ x[59];
  assign t[208] = t[251] ^ x[60];
  assign t[209] = t[252] ^ x[65];
  assign t[20] = t[12] ^ t[23];
  assign t[210] = t[253] ^ x[66];
  assign t[211] = t[254] ^ x[67];
  assign t[212] = t[255] ^ x[68];
  assign t[213] = t[256] ^ x[73];
  assign t[214] = t[257] ^ x[74];
  assign t[215] = t[258] ^ x[75];
  assign t[216] = t[259] ^ x[76];
  assign t[217] = t[260] ^ x[77];
  assign t[218] = t[261] ^ x[78];
  assign t[219] = t[262] ^ x[79];
  assign t[21] = x[7] ? t[28] : t[27];
  assign t[220] = t[263] ^ x[80];
  assign t[221] = t[264] ^ x[81];
  assign t[222] = t[265] ^ x[82];
  assign t[223] = t[266] ^ x[83];
  assign t[224] = t[267] ^ x[84];
  assign t[225] = t[268] ^ x[85];
  assign t[226] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[227] = (x[2]);
  assign t[228] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[229] = (x[11]);
  assign t[22] = x[7] ? t[30] : t[29];
  assign t[230] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[231] = (x[14]);
  assign t[232] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[233] = (x[17]);
  assign t[234] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[235] = (x[20]);
  assign t[236] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[237] = (x[24]);
  assign t[238] = (x[1]);
  assign t[239] = (x[26]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[240] = (x[23]);
  assign t[241] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[242] = (x[35]);
  assign t[243] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[244] = (x[43]);
  assign t[245] = (x[3]);
  assign t[246] = (x[0]);
  assign t[247] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[248] = (x[53]);
  assign t[249] = (x[25]);
  assign t[24] = t[33] ^ t[34];
  assign t[250] = (x[37]);
  assign t[251] = (x[34]);
  assign t[252] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[253] = (x[62]);
  assign t[254] = (x[45]);
  assign t[255] = (x[42]);
  assign t[256] = (x[69] & ~x[70] & ~x[71] & ~x[72]) | (~x[69] & x[70] & ~x[71] & ~x[72]) | (~x[69] & ~x[70] & x[71] & ~x[72]) | (~x[69] & ~x[70] & ~x[71] & x[72]) | (x[69] & x[70] & x[71] & ~x[72]) | (x[69] & x[70] & ~x[71] & x[72]) | (x[69] & ~x[70] & x[71] & x[72]) | (~x[69] & x[70] & x[71] & x[72]);
  assign t[257] = (x[70]);
  assign t[258] = (x[55]);
  assign t[259] = (x[52]);
  assign t[25] = ~(t[35] & t[36]);
  assign t[260] = (x[36]);
  assign t[261] = (x[64]);
  assign t[262] = (x[61]);
  assign t[263] = (x[44]);
  assign t[264] = (x[72]);
  assign t[265] = (x[69]);
  assign t[266] = (x[54]);
  assign t[267] = (x[63]);
  assign t[268] = (x[71]);
  assign t[26] = ~(t[37] & t[92]);
  assign t[27] = ~(t[38] & t[39]);
  assign t[28] = t[40] ^ t[41];
  assign t[29] = ~(t[42] & t[43]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[44] ^ t[45];
  assign t[31] = ~(t[46] & t[47]);
  assign t[32] = ~(t[48] & t[93]);
  assign t[33] = t[49] ? x[31] : x[30];
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = ~(t[94]);
  assign t[36] = ~(t[95]);
  assign t[37] = ~(t[52] & t[53]);
  assign t[38] = ~(t[54] & t[55]);
  assign t[39] = ~(t[56] & t[96]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[49] ? x[41] : x[40];
  assign t[41] = ~(t[57] & t[58]);
  assign t[42] = ~(t[59] & t[60]);
  assign t[43] = ~(t[61] & t[97]);
  assign t[44] = t[62] ? x[49] : x[48];
  assign t[45] = ~(t[63] & t[64]);
  assign t[46] = ~(t[98]);
  assign t[47] = ~(t[99]);
  assign t[48] = ~(t[65] & t[66]);
  assign t[49] = ~(t[67]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[68] & t[69]);
  assign t[51] = ~(t[70] & t[100]);
  assign t[52] = ~(t[95] & t[94]);
  assign t[53] = ~(t[101]);
  assign t[54] = ~(t[102]);
  assign t[55] = ~(t[103]);
  assign t[56] = ~(t[71] & t[72]);
  assign t[57] = ~(t[73] & t[74]);
  assign t[58] = ~(t[75] & t[104]);
  assign t[59] = ~(t[105]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[106]);
  assign t[61] = ~(t[76] & t[77]);
  assign t[62] = ~(t[67]);
  assign t[63] = ~(t[78] & t[79]);
  assign t[64] = ~(t[80] & t[107]);
  assign t[65] = ~(t[99] & t[98]);
  assign t[66] = ~(t[87]);
  assign t[67] = ~(t[88]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[109]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[81] & t[82]);
  assign t[71] = ~(t[103] & t[102]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[112]);
  assign t[75] = ~(t[83] & t[84]);
  assign t[76] = ~(t[106] & t[105]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[115]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[85] & t[86]);
  assign t[81] = ~(t[109] & t[108]);
  assign t[82] = ~(t[116]);
  assign t[83] = ~(t[112] & t[111]);
  assign t[84] = ~(t[117]);
  assign t[85] = ~(t[115] & t[114]);
  assign t[86] = ~(t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [79:0] x;
 output y;

 wire [225:0] t;
  assign t[0] = t[1] ? t[2] : t[74];
  assign t[100] = t[126] ^ x[5];
  assign t[101] = t[127] ^ x[13];
  assign t[102] = t[128] ^ x[16];
  assign t[103] = t[129] ^ x[19];
  assign t[104] = t[130] ^ x[22];
  assign t[105] = t[131] ^ x[28];
  assign t[106] = t[132] ^ x[29];
  assign t[107] = t[133] ^ x[30];
  assign t[108] = t[134] ^ x[31];
  assign t[109] = t[135] ^ x[34];
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[136] ^ x[40];
  assign t[111] = t[137] ^ x[41];
  assign t[112] = t[138] ^ x[49];
  assign t[113] = t[139] ^ x[50];
  assign t[114] = t[140] ^ x[53];
  assign t[115] = t[141] ^ x[59];
  assign t[116] = t[142] ^ x[60];
  assign t[117] = t[143] ^ x[61];
  assign t[118] = t[144] ^ x[67];
  assign t[119] = t[145] ^ x[68];
  assign t[11] = ~(x[6]);
  assign t[120] = t[146] ^ x[69];
  assign t[121] = t[147] ^ x[75];
  assign t[122] = t[148] ^ x[76];
  assign t[123] = t[149] ^ x[77];
  assign t[124] = t[150] ^ x[78];
  assign t[125] = t[151] ^ x[79];
  assign t[126] = (~t[152] & t[153]);
  assign t[127] = (~t[154] & t[155]);
  assign t[128] = (~t[156] & t[157]);
  assign t[129] = (~t[158] & t[159]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (~t[160] & t[161]);
  assign t[131] = (~t[162] & t[163]);
  assign t[132] = (~t[162] & t[164]);
  assign t[133] = (~t[152] & t[165]);
  assign t[134] = (~t[152] & t[166]);
  assign t[135] = (~t[162] & t[167]);
  assign t[136] = (~t[168] & t[169]);
  assign t[137] = (~t[168] & t[170]);
  assign t[138] = (~t[171] & t[172]);
  assign t[139] = (~t[171] & t[173]);
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = (~t[152] & t[174]);
  assign t[141] = (~t[175] & t[176]);
  assign t[142] = (~t[175] & t[177]);
  assign t[143] = (~t[168] & t[178]);
  assign t[144] = (~t[179] & t[180]);
  assign t[145] = (~t[179] & t[181]);
  assign t[146] = (~t[171] & t[182]);
  assign t[147] = (~t[183] & t[184]);
  assign t[148] = (~t[183] & t[185]);
  assign t[149] = (~t[175] & t[186]);
  assign t[14] = x[7] ? t[21] : t[20];
  assign t[150] = (~t[179] & t[187]);
  assign t[151] = (~t[183] & t[188]);
  assign t[152] = t[189] ^ x[4];
  assign t[153] = t[190] ^ x[5];
  assign t[154] = t[191] ^ x[12];
  assign t[155] = t[192] ^ x[13];
  assign t[156] = t[193] ^ x[15];
  assign t[157] = t[194] ^ x[16];
  assign t[158] = t[195] ^ x[18];
  assign t[159] = t[196] ^ x[19];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[197] ^ x[21];
  assign t[161] = t[198] ^ x[22];
  assign t[162] = t[199] ^ x[27];
  assign t[163] = t[200] ^ x[28];
  assign t[164] = t[201] ^ x[29];
  assign t[165] = t[202] ^ x[30];
  assign t[166] = t[203] ^ x[31];
  assign t[167] = t[204] ^ x[34];
  assign t[168] = t[205] ^ x[39];
  assign t[169] = t[206] ^ x[40];
  assign t[16] = ~(t[75] & t[76]);
  assign t[170] = t[207] ^ x[41];
  assign t[171] = t[208] ^ x[48];
  assign t[172] = t[209] ^ x[49];
  assign t[173] = t[210] ^ x[50];
  assign t[174] = t[211] ^ x[53];
  assign t[175] = t[212] ^ x[58];
  assign t[176] = t[213] ^ x[59];
  assign t[177] = t[214] ^ x[60];
  assign t[178] = t[215] ^ x[61];
  assign t[179] = t[216] ^ x[66];
  assign t[17] = ~(t[77] & t[78]);
  assign t[180] = t[217] ^ x[67];
  assign t[181] = t[218] ^ x[68];
  assign t[182] = t[219] ^ x[69];
  assign t[183] = t[220] ^ x[74];
  assign t[184] = t[221] ^ x[75];
  assign t[185] = t[222] ^ x[76];
  assign t[186] = t[223] ^ x[77];
  assign t[187] = t[224] ^ x[78];
  assign t[188] = t[225] ^ x[79];
  assign t[189] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[1]);
  assign t[191] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[192] = (x[11]);
  assign t[193] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[194] = (x[14]);
  assign t[195] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[196] = (x[17]);
  assign t[197] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[198] = (x[20]);
  assign t[199] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[19] = x[7] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = (x[25]);
  assign t[201] = (x[23]);
  assign t[202] = (x[2]);
  assign t[203] = (x[0]);
  assign t[204] = (x[26]);
  assign t[205] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[206] = (x[37]);
  assign t[207] = (x[35]);
  assign t[208] = (x[44] & ~x[45] & ~x[46] & ~x[47]) | (~x[44] & x[45] & ~x[46] & ~x[47]) | (~x[44] & ~x[45] & x[46] & ~x[47]) | (~x[44] & ~x[45] & ~x[46] & x[47]) | (x[44] & x[45] & x[46] & ~x[47]) | (x[44] & x[45] & ~x[46] & x[47]) | (x[44] & ~x[45] & x[46] & x[47]) | (~x[44] & x[45] & x[46] & x[47]);
  assign t[209] = (x[46]);
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = (x[44]);
  assign t[211] = (x[3]);
  assign t[212] = (x[54] & ~x[55] & ~x[56] & ~x[57]) | (~x[54] & x[55] & ~x[56] & ~x[57]) | (~x[54] & ~x[55] & x[56] & ~x[57]) | (~x[54] & ~x[55] & ~x[56] & x[57]) | (x[54] & x[55] & x[56] & ~x[57]) | (x[54] & x[55] & ~x[56] & x[57]) | (x[54] & ~x[55] & x[56] & x[57]) | (~x[54] & x[55] & x[56] & x[57]);
  assign t[213] = (x[56]);
  assign t[214] = (x[54]);
  assign t[215] = (x[38]);
  assign t[216] = (x[62] & ~x[63] & ~x[64] & ~x[65]) | (~x[62] & x[63] & ~x[64] & ~x[65]) | (~x[62] & ~x[63] & x[64] & ~x[65]) | (~x[62] & ~x[63] & ~x[64] & x[65]) | (x[62] & x[63] & x[64] & ~x[65]) | (x[62] & x[63] & ~x[64] & x[65]) | (x[62] & ~x[63] & x[64] & x[65]) | (~x[62] & x[63] & x[64] & x[65]);
  assign t[217] = (x[64]);
  assign t[218] = (x[62]);
  assign t[219] = (x[47]);
  assign t[21] = t[12] ^ t[25];
  assign t[220] = (x[70] & ~x[71] & ~x[72] & ~x[73]) | (~x[70] & x[71] & ~x[72] & ~x[73]) | (~x[70] & ~x[71] & x[72] & ~x[73]) | (~x[70] & ~x[71] & ~x[72] & x[73]) | (x[70] & x[71] & x[72] & ~x[73]) | (x[70] & x[71] & ~x[72] & x[73]) | (x[70] & ~x[71] & x[72] & x[73]) | (~x[70] & x[71] & x[72] & x[73]);
  assign t[221] = (x[72]);
  assign t[222] = (x[70]);
  assign t[223] = (x[57]);
  assign t[224] = (x[65]);
  assign t[225] = (x[73]);
  assign t[22] = x[7] ? t[30] : t[29];
  assign t[23] = x[7] ? t[32] : t[31];
  assign t[24] = ~(t[77]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[79] & t[37]);
  assign t[28] = ~(t[80] & t[38]);
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[43] & t[44]);
  assign t[32] = t[45] ^ t[46];
  assign t[33] = ~(t[81] & t[47]);
  assign t[34] = ~(t[82] & t[48]);
  assign t[35] = t[49] ? x[33] : x[32];
  assign t[36] = ~(t[50] & t[51]);
  assign t[37] = ~(t[83]);
  assign t[38] = ~(t[83] & t[52]);
  assign t[39] = ~(t[84] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[85] & t[54]);
  assign t[41] = t[55] ? x[43] : x[42];
  assign t[42] = ~(t[56] & t[57]);
  assign t[43] = ~(t[86] & t[58]);
  assign t[44] = ~(t[87] & t[59]);
  assign t[45] = t[49] ? x[52] : x[51];
  assign t[46] = ~(t[60] & t[61]);
  assign t[47] = ~(t[88]);
  assign t[48] = ~(t[88] & t[62]);
  assign t[49] = ~(t[24]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[89] & t[63]);
  assign t[51] = ~(t[90] & t[64]);
  assign t[52] = ~(t[79]);
  assign t[53] = ~(t[91]);
  assign t[54] = ~(t[91] & t[65]);
  assign t[55] = ~(t[24]);
  assign t[56] = ~(t[92] & t[66]);
  assign t[57] = ~(t[93] & t[67]);
  assign t[58] = ~(t[94]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[95] & t[69]);
  assign t[61] = ~(t[96] & t[70]);
  assign t[62] = ~(t[81]);
  assign t[63] = ~(t[97]);
  assign t[64] = ~(t[97] & t[71]);
  assign t[65] = ~(t[84]);
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[98] & t[72]);
  assign t[68] = ~(t[86]);
  assign t[69] = ~(t[99]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[99] & t[73]);
  assign t[71] = ~(t[89]);
  assign t[72] = ~(t[92]);
  assign t[73] = ~(t[95]);
  assign t[74] = (t[100]);
  assign t[75] = (t[101]);
  assign t[76] = (t[102]);
  assign t[77] = (t[103]);
  assign t[78] = (t[104]);
  assign t[79] = (t[105]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[106]);
  assign t[81] = (t[107]);
  assign t[82] = (t[108]);
  assign t[83] = (t[109]);
  assign t[84] = (t[110]);
  assign t[85] = (t[111]);
  assign t[86] = (t[112]);
  assign t[87] = (t[113]);
  assign t[88] = (t[114]);
  assign t[89] = (t[115]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[116]);
  assign t[91] = (t[117]);
  assign t[92] = (t[118]);
  assign t[93] = (t[119]);
  assign t[94] = (t[120]);
  assign t[95] = (t[121]);
  assign t[96] = (t[122]);
  assign t[97] = (t[123]);
  assign t[98] = (t[124]);
  assign t[99] = (t[125]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [85:0] x;
 output y;

 wire [343:0] t;
  assign t[0] = t[1] ? t[2] : t[162];
  assign t[100] = t[63] & t[163];
  assign t[101] = ~(t[185]);
  assign t[102] = ~(t[177] | t[178]);
  assign t[103] = ~(t[186]);
  assign t[104] = ~(t[187]);
  assign t[105] = ~(t[126] | t[127]);
  assign t[106] = ~(t[43] | t[128]);
  assign t[107] = ~(t[42] | t[129]);
  assign t[108] = ~(t[188]);
  assign t[109] = ~(t[180] | t[181]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[189]);
  assign t[111] = ~(t[190]);
  assign t[112] = ~(t[130] | t[131]);
  assign t[113] = ~(t[132] | t[133]);
  assign t[114] = ~(t[117] | t[134]);
  assign t[115] = ~(t[191]);
  assign t[116] = ~(t[183] | t[184]);
  assign t[117] = ~(t[63] | t[135]);
  assign t[118] = ~(t[63] | t[136]);
  assign t[119] = t[44] | t[137];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[138] & t[139]);
  assign t[121] = x[7] & t[164];
  assign t[122] = ~(x[7] | t[164]);
  assign t[123] = ~(t[166]);
  assign t[124] = t[163] ? t[95] : t[94];
  assign t[125] = t[163] ? t[141] : t[140];
  assign t[126] = ~(t[192]);
  assign t[127] = ~(t[186] | t[187]);
  assign t[128] = ~(t[63] | t[142]);
  assign t[129] = ~(t[114] & t[139]);
  assign t[12] = ~(t[18] ^ t[15]);
  assign t[130] = ~(t[193]);
  assign t[131] = ~(t[189] | t[190]);
  assign t[132] = ~(t[106] & t[143]);
  assign t[133] = ~(t[144] & t[139]);
  assign t[134] = ~(t[63] | t[145]);
  assign t[135] = t[163] ? t[93] : t[94];
  assign t[136] = t[163] ? t[140] : t[146];
  assign t[137] = ~(t[63] | t[147]);
  assign t[138] = ~(t[148] | t[149]);
  assign t[139] = t[66] | t[150];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = ~(x[7] & t[151]);
  assign t[141] = ~(t[152] & t[123]);
  assign t[142] = t[163] ? t[141] : t[153];
  assign t[143] = ~(t[66] & t[154]);
  assign t[144] = ~(t[155] & t[156]);
  assign t[145] = t[163] ? t[95] : t[96];
  assign t[146] = ~(t[166] & t[152]);
  assign t[147] = t[163] ? t[146] : t[140];
  assign t[148] = ~(t[157]);
  assign t[149] = ~(t[63] | t[158]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[163] ? t[140] : t[141];
  assign t[151] = ~(t[164] | t[166]);
  assign t[152] = ~(x[7] | t[159]);
  assign t[153] = ~(x[7] & t[99]);
  assign t[154] = ~(t[140] & t[146]);
  assign t[155] = t[166] & t[160];
  assign t[156] = t[122] | t[121];
  assign t[157] = ~(t[160] & t[161]);
  assign t[158] = t[163] ? t[153] : t[141];
  assign t[159] = ~(t[164]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = ~(t[66] | t[163]);
  assign t[161] = ~(t[146] & t[153]);
  assign t[162] = (t[194]);
  assign t[163] = (t[195]);
  assign t[164] = (t[196]);
  assign t[165] = (t[197]);
  assign t[166] = (t[198]);
  assign t[167] = (t[199]);
  assign t[168] = (t[200]);
  assign t[169] = (t[201]);
  assign t[16] = ~(t[163] & t[164]);
  assign t[170] = (t[202]);
  assign t[171] = (t[203]);
  assign t[172] = (t[204]);
  assign t[173] = (t[205]);
  assign t[174] = (t[206]);
  assign t[175] = (t[207]);
  assign t[176] = (t[208]);
  assign t[177] = (t[209]);
  assign t[178] = (t[210]);
  assign t[179] = (t[211]);
  assign t[17] = ~(t[165] & t[166]);
  assign t[180] = (t[212]);
  assign t[181] = (t[213]);
  assign t[182] = (t[214]);
  assign t[183] = (t[215]);
  assign t[184] = (t[216]);
  assign t[185] = (t[217]);
  assign t[186] = (t[218]);
  assign t[187] = (t[219]);
  assign t[188] = (t[220]);
  assign t[189] = (t[221]);
  assign t[18] = x[7] ? t[26] : t[25];
  assign t[190] = (t[222]);
  assign t[191] = (t[223]);
  assign t[192] = (t[224]);
  assign t[193] = (t[225]);
  assign t[194] = t[226] ^ x[5];
  assign t[195] = t[227] ^ x[13];
  assign t[196] = t[228] ^ x[16];
  assign t[197] = t[229] ^ x[19];
  assign t[198] = t[230] ^ x[22];
  assign t[199] = t[231] ^ x[28];
  assign t[19] = t[27] ? x[9] : x[10];
  assign t[1] = ~(t[3]);
  assign t[200] = t[232] ^ x[29];
  assign t[201] = t[233] ^ x[30];
  assign t[202] = t[234] ^ x[31];
  assign t[203] = t[235] ^ x[37];
  assign t[204] = t[236] ^ x[43];
  assign t[205] = t[237] ^ x[44];
  assign t[206] = t[238] ^ x[45];
  assign t[207] = t[239] ^ x[51];
  assign t[208] = t[240] ^ x[54];
  assign t[209] = t[241] ^ x[55];
  assign t[20] = ~(t[28] & t[29]);
  assign t[210] = t[242] ^ x[56];
  assign t[211] = t[243] ^ x[62];
  assign t[212] = t[244] ^ x[65];
  assign t[213] = t[245] ^ x[66];
  assign t[214] = t[246] ^ x[72];
  assign t[215] = t[247] ^ x[75];
  assign t[216] = t[248] ^ x[76];
  assign t[217] = t[249] ^ x[77];
  assign t[218] = t[250] ^ x[78];
  assign t[219] = t[251] ^ x[79];
  assign t[21] = ~(t[30] | t[31]);
  assign t[220] = t[252] ^ x[80];
  assign t[221] = t[253] ^ x[81];
  assign t[222] = t[254] ^ x[82];
  assign t[223] = t[255] ^ x[83];
  assign t[224] = t[256] ^ x[84];
  assign t[225] = t[257] ^ x[85];
  assign t[226] = (~t[258] & t[259]);
  assign t[227] = (~t[260] & t[261]);
  assign t[228] = (~t[262] & t[263]);
  assign t[229] = (~t[264] & t[265]);
  assign t[22] = ~(t[25] ^ t[13]);
  assign t[230] = (~t[266] & t[267]);
  assign t[231] = (~t[268] & t[269]);
  assign t[232] = (~t[258] & t[270]);
  assign t[233] = (~t[268] & t[271]);
  assign t[234] = (~t[268] & t[272]);
  assign t[235] = (~t[273] & t[274]);
  assign t[236] = (~t[275] & t[276]);
  assign t[237] = (~t[258] & t[277]);
  assign t[238] = (~t[258] & t[278]);
  assign t[239] = (~t[279] & t[280]);
  assign t[23] = x[7] ? t[33] : t[32];
  assign t[240] = (~t[268] & t[281]);
  assign t[241] = (~t[273] & t[282]);
  assign t[242] = (~t[273] & t[283]);
  assign t[243] = (~t[284] & t[285]);
  assign t[244] = (~t[275] & t[286]);
  assign t[245] = (~t[275] & t[287]);
  assign t[246] = (~t[288] & t[289]);
  assign t[247] = (~t[279] & t[290]);
  assign t[248] = (~t[279] & t[291]);
  assign t[249] = (~t[273] & t[292]);
  assign t[24] = x[7] ? t[35] : t[34];
  assign t[250] = (~t[284] & t[293]);
  assign t[251] = (~t[284] & t[294]);
  assign t[252] = (~t[275] & t[295]);
  assign t[253] = (~t[288] & t[296]);
  assign t[254] = (~t[288] & t[297]);
  assign t[255] = (~t[279] & t[298]);
  assign t[256] = (~t[284] & t[299]);
  assign t[257] = (~t[288] & t[300]);
  assign t[258] = t[301] ^ x[4];
  assign t[259] = t[302] ^ x[5];
  assign t[25] = ~(t[36] | t[37]);
  assign t[260] = t[303] ^ x[12];
  assign t[261] = t[304] ^ x[13];
  assign t[262] = t[305] ^ x[15];
  assign t[263] = t[306] ^ x[16];
  assign t[264] = t[307] ^ x[18];
  assign t[265] = t[308] ^ x[19];
  assign t[266] = t[309] ^ x[21];
  assign t[267] = t[310] ^ x[22];
  assign t[268] = t[311] ^ x[27];
  assign t[269] = t[312] ^ x[28];
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = t[313] ^ x[29];
  assign t[271] = t[314] ^ x[30];
  assign t[272] = t[315] ^ x[31];
  assign t[273] = t[316] ^ x[36];
  assign t[274] = t[317] ^ x[37];
  assign t[275] = t[318] ^ x[42];
  assign t[276] = t[319] ^ x[43];
  assign t[277] = t[320] ^ x[44];
  assign t[278] = t[321] ^ x[45];
  assign t[279] = t[322] ^ x[50];
  assign t[27] = ~(t[40]);
  assign t[280] = t[323] ^ x[51];
  assign t[281] = t[324] ^ x[54];
  assign t[282] = t[325] ^ x[55];
  assign t[283] = t[326] ^ x[56];
  assign t[284] = t[327] ^ x[61];
  assign t[285] = t[328] ^ x[62];
  assign t[286] = t[329] ^ x[65];
  assign t[287] = t[330] ^ x[66];
  assign t[288] = t[331] ^ x[71];
  assign t[289] = t[332] ^ x[72];
  assign t[28] = ~(t[41] | t[42]);
  assign t[290] = t[333] ^ x[75];
  assign t[291] = t[334] ^ x[76];
  assign t[292] = t[335] ^ x[77];
  assign t[293] = t[336] ^ x[78];
  assign t[294] = t[337] ^ x[79];
  assign t[295] = t[338] ^ x[80];
  assign t[296] = t[339] ^ x[81];
  assign t[297] = t[340] ^ x[82];
  assign t[298] = t[341] ^ x[83];
  assign t[299] = t[342] ^ x[84];
  assign t[29] = ~(t[43] | t[44]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[343] ^ x[85];
  assign t[301] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[302] = (x[0]);
  assign t[303] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[304] = (x[11]);
  assign t[305] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[306] = (x[14]);
  assign t[307] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[308] = (x[17]);
  assign t[309] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[30] = ~(t[45] | t[46]);
  assign t[310] = (x[20]);
  assign t[311] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[312] = (x[24]);
  assign t[313] = (x[1]);
  assign t[314] = (x[25]);
  assign t[315] = (x[26]);
  assign t[316] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[317] = (x[33]);
  assign t[318] = (x[38] & ~x[39] & ~x[40] & ~x[41]) | (~x[38] & x[39] & ~x[40] & ~x[41]) | (~x[38] & ~x[39] & x[40] & ~x[41]) | (~x[38] & ~x[39] & ~x[40] & x[41]) | (x[38] & x[39] & x[40] & ~x[41]) | (x[38] & x[39] & ~x[40] & x[41]) | (x[38] & ~x[39] & x[40] & x[41]) | (~x[38] & x[39] & x[40] & x[41]);
  assign t[319] = (x[39]);
  assign t[31] = ~(t[167] | t[47]);
  assign t[320] = (x[2]);
  assign t[321] = (x[3]);
  assign t[322] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[323] = (x[47]);
  assign t[324] = (x[23]);
  assign t[325] = (x[34]);
  assign t[326] = (x[35]);
  assign t[327] = (x[57] & ~x[58] & ~x[59] & ~x[60]) | (~x[57] & x[58] & ~x[59] & ~x[60]) | (~x[57] & ~x[58] & x[59] & ~x[60]) | (~x[57] & ~x[58] & ~x[59] & x[60]) | (x[57] & x[58] & x[59] & ~x[60]) | (x[57] & x[58] & ~x[59] & x[60]) | (x[57] & ~x[58] & x[59] & x[60]) | (~x[57] & x[58] & x[59] & x[60]);
  assign t[328] = (x[58]);
  assign t[329] = (x[40]);
  assign t[32] = ~(t[48] | t[49]);
  assign t[330] = (x[41]);
  assign t[331] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[332] = (x[68]);
  assign t[333] = (x[48]);
  assign t[334] = (x[49]);
  assign t[335] = (x[32]);
  assign t[336] = (x[59]);
  assign t[337] = (x[60]);
  assign t[338] = (x[38]);
  assign t[339] = (x[69]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[340] = (x[70]);
  assign t[341] = (x[46]);
  assign t[342] = (x[57]);
  assign t[343] = (x[67]);
  assign t[34] = ~(t[52] | t[53]);
  assign t[35] = ~(t[54] ^ t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = ~(t[168] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = ~(t[61] ^ t[62]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[165]);
  assign t[41] = ~(t[63] | t[64]);
  assign t[42] = ~(t[63] | t[65]);
  assign t[43] = ~(t[66] | t[67]);
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = ~(t[169]);
  assign t[46] = ~(t[170]);
  assign t[47] = ~(t[70] | t[71]);
  assign t[48] = ~(t[72] | t[73]);
  assign t[49] = ~(t[171] | t[74]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[75] | t[76]);
  assign t[51] = ~(t[77] ^ t[78]);
  assign t[52] = ~(t[79] | t[80]);
  assign t[53] = ~(t[172] | t[81]);
  assign t[54] = ~(t[82] | t[83]);
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = ~(t[173]);
  assign t[57] = ~(t[174]);
  assign t[58] = ~(t[86] | t[87]);
  assign t[59] = ~(t[88] | t[89]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[175] | t[90]);
  assign t[61] = t[27] ? x[53] : x[52];
  assign t[62] = ~(t[91] & t[92]);
  assign t[63] = ~(t[66]);
  assign t[64] = t[163] ? t[94] : t[93];
  assign t[65] = t[163] ? t[96] : t[95];
  assign t[66] = ~(t[165]);
  assign t[67] = t[163] ? t[94] : t[95];
  assign t[68] = ~(t[97] | t[98]);
  assign t[69] = ~(t[99] & t[100]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[176]);
  assign t[71] = ~(t[169] | t[170]);
  assign t[72] = ~(t[177]);
  assign t[73] = ~(t[178]);
  assign t[74] = ~(t[101] | t[102]);
  assign t[75] = ~(t[103] | t[104]);
  assign t[76] = ~(t[179] | t[105]);
  assign t[77] = t[27] ? x[64] : x[63];
  assign t[78] = ~(t[106] & t[107]);
  assign t[79] = ~(t[180]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[181]);
  assign t[81] = ~(t[108] | t[109]);
  assign t[82] = ~(t[110] | t[111]);
  assign t[83] = ~(t[182] | t[112]);
  assign t[84] = t[27] ? x[74] : x[73];
  assign t[85] = ~(t[113] & t[114]);
  assign t[86] = ~(t[162]);
  assign t[87] = ~(t[173] | t[174]);
  assign t[88] = ~(t[183]);
  assign t[89] = ~(t[184]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[115] | t[116]);
  assign t[91] = ~(t[117] | t[118]);
  assign t[92] = ~(t[119] | t[120]);
  assign t[93] = ~(t[121] & t[166]);
  assign t[94] = ~(t[122] & t[123]);
  assign t[95] = ~(t[121] & t[123]);
  assign t[96] = ~(t[122] & t[166]);
  assign t[97] = ~(t[66] | t[124]);
  assign t[98] = ~(t[66] | t[125]);
  assign t[99] = ~(t[164] | t[123]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [172:0] x;
 output y;

 wire [679:0] t;
  assign t[0] = t[1] ? t[2] : t[410];
  assign t[100] = ~(t[147] & t[148]);
  assign t[101] = ~(t[432]);
  assign t[102] = ~(t[433]);
  assign t[103] = ~(t[149] | t[150]);
  assign t[104] = t[413] ? x[89] : x[88];
  assign t[105] = t[151] | t[152];
  assign t[106] = ~(t[434]);
  assign t[107] = ~(t[422] | t[423]);
  assign t[108] = ~(t[435]);
  assign t[109] = ~(t[436]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[153] | t[154]);
  assign t[111] = ~(t[140] | t[155]);
  assign t[112] = ~(t[156] | t[85]);
  assign t[113] = ~(t[437]);
  assign t[114] = ~(t[438]);
  assign t[115] = ~(t[157] | t[158]);
  assign t[116] = ~(t[159] | t[160]);
  assign t[117] = ~(t[439] | t[161]);
  assign t[118] = t[30] ? x[102] : x[101];
  assign t[119] = ~(t[162] & t[163]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[440]);
  assign t[121] = ~(t[441]);
  assign t[122] = ~(t[164] | t[165]);
  assign t[123] = ~(t[166] | t[167]);
  assign t[124] = ~(t[442] | t[168]);
  assign t[125] = t[30] ? x[112] : x[111];
  assign t[126] = ~(t[169] & t[170]);
  assign t[127] = ~(t[413]);
  assign t[128] = ~(t[171] & t[172]);
  assign t[129] = ~(t[173] & t[414]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[414] & t[174]);
  assign t[131] = ~(x[7] & t[175]);
  assign t[132] = ~(t[176] | t[142]);
  assign t[133] = ~(t[177] & t[178]);
  assign t[134] = t[411] ? t[130] : t[131];
  assign t[135] = ~(t[179]);
  assign t[136] = ~(t[82] | t[180]);
  assign t[137] = t[411] ? t[131] : t[181];
  assign t[138] = ~(t[443]);
  assign t[139] = ~(t[428] | t[429]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[82] | t[182]);
  assign t[141] = ~(t[31] & t[183]);
  assign t[142] = ~(t[127] | t[184]);
  assign t[143] = t[155] | t[135];
  assign t[144] = ~(t[444]);
  assign t[145] = ~(t[430] | t[431]);
  assign t[146] = ~(t[49]);
  assign t[147] = ~(t[151] | t[185]);
  assign t[148] = ~(t[140]);
  assign t[149] = ~(t[445]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[432] | t[433]);
  assign t[151] = ~(t[179] & t[133]);
  assign t[152] = ~(t[111] & t[186]);
  assign t[153] = ~(t[446]);
  assign t[154] = ~(t[435] | t[436]);
  assign t[155] = ~(t[82] | t[187]);
  assign t[156] = ~(t[127] | t[188]);
  assign t[157] = ~(t[447]);
  assign t[158] = ~(t[437] | t[438]);
  assign t[159] = ~(t[448]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[449]);
  assign t[161] = ~(t[189] | t[190]);
  assign t[162] = ~(t[156] | t[191]);
  assign t[163] = ~(t[155] | t[192]);
  assign t[164] = ~(t[450]);
  assign t[165] = ~(t[440] | t[441]);
  assign t[166] = ~(t[451]);
  assign t[167] = ~(t[452]);
  assign t[168] = ~(t[193] | t[194]);
  assign t[169] = ~(t[195] | t[196]);
  assign t[16] = ~(t[411] & t[412]);
  assign t[170] = ~(t[50] | t[197]);
  assign t[171] = ~(x[7] | t[412]);
  assign t[172] = ~(t[414]);
  assign t[173] = x[7] & t[412];
  assign t[174] = ~(x[7] | t[198]);
  assign t[175] = ~(t[412] | t[414]);
  assign t[176] = ~(t[127] | t[199]);
  assign t[177] = ~(t[412] | t[172]);
  assign t[178] = t[82] & t[411];
  assign t[179] = ~(t[200] & t[201]);
  assign t[17] = ~(t[413] & t[414]);
  assign t[180] = t[411] ? t[202] : t[181];
  assign t[181] = ~(t[174] & t[172]);
  assign t[182] = t[411] ? t[128] : t[129];
  assign t[183] = ~(t[203] & t[204]);
  assign t[184] = t[411] ? t[181] : t[131];
  assign t[185] = ~(t[205] & t[88]);
  assign t[186] = ~(t[51] | t[197]);
  assign t[187] = t[411] ? t[207] : t[206];
  assign t[188] = t[411] ? t[128] : t[206];
  assign t[189] = ~(t[453]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[448] | t[449]);
  assign t[191] = ~(t[82] | t[208]);
  assign t[192] = ~(t[170] & t[88]);
  assign t[193] = ~(t[454]);
  assign t[194] = ~(t[451] | t[452]);
  assign t[195] = ~(t[162] & t[209]);
  assign t[196] = ~(t[183] & t[88]);
  assign t[197] = ~(t[82] | t[210]);
  assign t[198] = ~(t[412]);
  assign t[199] = t[411] ? t[206] : t[128];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[127] | t[411]);
  assign t[201] = ~(t[130] & t[202]);
  assign t[202] = ~(x[7] & t[177]);
  assign t[203] = t[414] & t[200];
  assign t[204] = t[171] | t[173];
  assign t[205] = ~(t[142]);
  assign t[206] = ~(t[173] & t[172]);
  assign t[207] = ~(t[171] & t[414]);
  assign t[208] = t[411] ? t[181] : t[202];
  assign t[209] = ~(t[127] & t[211]);
  assign t[20] = t[30] ? x[9] : x[10];
  assign t[210] = t[411] ? t[206] : t[207];
  assign t[211] = ~(t[131] & t[130]);
  assign t[212] = t[1] ? t[213] : t[455];
  assign t[213] = x[6] ? t[215] : t[214];
  assign t[214] = x[7] ? t[217] : t[216];
  assign t[215] = t[218] ^ x[126];
  assign t[216] = t[219] ^ t[220];
  assign t[217] = ~(t[221] ^ t[222]);
  assign t[218] = x[127] ^ x[128];
  assign t[219] = t[30] ? x[127] : x[128];
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = ~(t[223] ^ t[224]);
  assign t[221] = x[7] ? t[226] : t[225];
  assign t[222] = ~(t[227] ^ t[228]);
  assign t[223] = x[7] ? t[230] : t[229];
  assign t[224] = ~(t[231] ^ t[232]);
  assign t[225] = ~(t[233] & t[234]);
  assign t[226] = t[235] ^ t[236];
  assign t[227] = x[7] ? t[238] : t[237];
  assign t[228] = x[7] ? t[240] : t[239];
  assign t[229] = ~(t[241] & t[242]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = t[243] ^ t[244];
  assign t[231] = x[7] ? t[246] : t[245];
  assign t[232] = x[7] ? t[248] : t[247];
  assign t[233] = ~(t[417] & t[55]);
  assign t[234] = ~(t[427] & t[249]);
  assign t[235] = t[250] ? x[130] : x[129];
  assign t[236] = ~(t[251] & t[252]);
  assign t[237] = ~(t[253] & t[254]);
  assign t[238] = t[255] ^ t[237];
  assign t[239] = ~(t[256] & t[257]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = t[258] ^ t[247];
  assign t[241] = ~(t[422] & t[68]);
  assign t[242] = ~(t[434] & t[259]);
  assign t[243] = t[146] ? x[132] : x[131];
  assign t[244] = ~(t[260] & t[261]);
  assign t[245] = ~(t[262] & t[263]);
  assign t[246] = t[264] ^ t[265];
  assign t[247] = ~(t[266] & t[267]);
  assign t[248] = t[268] ^ t[269];
  assign t[249] = ~(t[418] & t[54]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = ~(t[49]);
  assign t[251] = ~(t[428] & t[92]);
  assign t[252] = ~(t[443] & t[270]);
  assign t[253] = ~(t[432] & t[102]);
  assign t[254] = ~(t[445] & t[271]);
  assign t[255] = t[413] ? x[134] : x[133];
  assign t[256] = ~(t[430] & t[97]);
  assign t[257] = ~(t[444] & t[272]);
  assign t[258] = t[413] ? x[136] : x[135];
  assign t[259] = ~(t[423] & t[67]);
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = ~(t[435] & t[109]);
  assign t[261] = ~(t[446] & t[273]);
  assign t[262] = ~(t[440] & t[121]);
  assign t[263] = ~(t[450] & t[274]);
  assign t[264] = t[250] ? x[138] : x[137];
  assign t[265] = ~(t[275] & t[276]);
  assign t[266] = ~(t[437] & t[114]);
  assign t[267] = ~(t[447] & t[277]);
  assign t[268] = t[30] ? x[140] : x[139];
  assign t[269] = ~(t[278] & t[279]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = ~(t[429] & t[91]);
  assign t[271] = ~(t[433] & t[101]);
  assign t[272] = ~(t[431] & t[96]);
  assign t[273] = ~(t[436] & t[108]);
  assign t[274] = ~(t[441] & t[120]);
  assign t[275] = ~(t[451] & t[167]);
  assign t[276] = ~(t[454] & t[280]);
  assign t[277] = ~(t[438] & t[113]);
  assign t[278] = ~(t[448] & t[160]);
  assign t[279] = ~(t[453] & t[281]);
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = ~(t[452] & t[166]);
  assign t[281] = ~(t[449] & t[159]);
  assign t[282] = t[1] ? t[283] : t[456];
  assign t[283] = x[6] ? t[285] : t[284];
  assign t[284] = x[7] ? t[287] : t[286];
  assign t[285] = t[288] ^ x[142];
  assign t[286] = t[289] ^ t[290];
  assign t[287] = ~(t[291] ^ t[292]);
  assign t[288] = x[143] ^ x[144];
  assign t[289] = t[30] ? x[143] : x[144];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = ~(t[293] ^ t[294]);
  assign t[291] = x[7] ? t[296] : t[295];
  assign t[292] = ~(t[297] ^ t[298]);
  assign t[293] = x[7] ? t[300] : t[299];
  assign t[294] = ~(t[301] ^ t[302]);
  assign t[295] = ~(t[303] & t[304]);
  assign t[296] = t[305] ^ t[306];
  assign t[297] = x[7] ? t[308] : t[307];
  assign t[298] = x[7] ? t[310] : t[309];
  assign t[299] = ~(t[311] & t[312]);
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[313] ^ t[314];
  assign t[301] = x[7] ? t[316] : t[315];
  assign t[302] = x[7] ? t[318] : t[317];
  assign t[303] = ~(t[55] & t[89]);
  assign t[304] = ~(t[319] & t[415]);
  assign t[305] = t[30] ? x[146] : x[145];
  assign t[306] = ~(t[320] & t[321]);
  assign t[307] = ~(t[322] & t[323]);
  assign t[308] = t[324] ^ t[317];
  assign t[309] = ~(t[325] & t[326]);
  assign t[30] = ~(t[49]);
  assign t[310] = t[327] ^ t[309];
  assign t[311] = ~(t[68] & t[106]);
  assign t[312] = ~(t[328] & t[416]);
  assign t[313] = t[413] ? x[148] : x[147];
  assign t[314] = ~(t[329] & t[330]);
  assign t[315] = ~(t[331] & t[332]);
  assign t[316] = t[333] ^ t[334];
  assign t[317] = ~(t[335] & t[336]);
  assign t[318] = t[337] ^ t[338];
  assign t[319] = ~(t[339] & t[54]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = ~(t[92] & t[138]);
  assign t[321] = ~(t[340] & t[419]);
  assign t[322] = ~(t[97] & t[144]);
  assign t[323] = ~(t[341] & t[420]);
  assign t[324] = t[413] ? x[150] : x[149];
  assign t[325] = ~(t[102] & t[149]);
  assign t[326] = ~(t[342] & t[421]);
  assign t[327] = t[413] ? x[152] : x[151];
  assign t[328] = ~(t[343] & t[67]);
  assign t[329] = ~(t[109] & t[153]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = ~(t[344] & t[424]);
  assign t[331] = ~(t[121] & t[164]);
  assign t[332] = ~(t[345] & t[426]);
  assign t[333] = t[30] ? x[154] : x[153];
  assign t[334] = ~(t[346] & t[347]);
  assign t[335] = ~(t[114] & t[157]);
  assign t[336] = ~(t[348] & t[425]);
  assign t[337] = t[146] ? x[156] : x[155];
  assign t[338] = ~(t[349] & t[350]);
  assign t[339] = ~(t[427] & t[418]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = ~(t[351] & t[91]);
  assign t[341] = ~(t[352] & t[96]);
  assign t[342] = ~(t[353] & t[101]);
  assign t[343] = ~(t[434] & t[423]);
  assign t[344] = ~(t[354] & t[108]);
  assign t[345] = ~(t[355] & t[120]);
  assign t[346] = ~(t[167] & t[193]);
  assign t[347] = ~(t[356] & t[442]);
  assign t[348] = ~(t[357] & t[113]);
  assign t[349] = ~(t[160] & t[189]);
  assign t[34] = ~(t[415] | t[56]);
  assign t[350] = ~(t[358] & t[439]);
  assign t[351] = ~(t[443] & t[429]);
  assign t[352] = ~(t[444] & t[431]);
  assign t[353] = ~(t[445] & t[433]);
  assign t[354] = ~(t[446] & t[436]);
  assign t[355] = ~(t[450] & t[441]);
  assign t[356] = ~(t[359] & t[166]);
  assign t[357] = ~(t[447] & t[438]);
  assign t[358] = ~(t[360] & t[159]);
  assign t[359] = ~(t[454] & t[452]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = ~(t[453] & t[449]);
  assign t[361] = t[1] ? t[362] : t[457];
  assign t[362] = x[6] ? t[364] : t[363];
  assign t[363] = x[7] ? t[366] : t[365];
  assign t[364] = t[367] ^ x[158];
  assign t[365] = t[368] ^ t[369];
  assign t[366] = ~(t[370] ^ t[371]);
  assign t[367] = x[159] ^ x[160];
  assign t[368] = t[30] ? x[159] : x[160];
  assign t[369] = ~(t[372] ^ t[373]);
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = x[7] ? t[375] : t[374];
  assign t[371] = ~(t[376] ^ t[377]);
  assign t[372] = x[7] ? t[379] : t[378];
  assign t[373] = ~(t[380] ^ t[381]);
  assign t[374] = ~(t[303] & t[382]);
  assign t[375] = t[383] ^ t[384];
  assign t[376] = x[7] ? t[386] : t[385];
  assign t[377] = x[7] ? t[388] : t[387];
  assign t[378] = ~(t[311] & t[389]);
  assign t[379] = t[390] ^ t[391];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = x[7] ? t[393] : t[392];
  assign t[381] = x[7] ? t[395] : t[394];
  assign t[382] = t[33] | t[415];
  assign t[383] = t[146] ? x[162] : x[161];
  assign t[384] = ~(t[320] & t[396]);
  assign t[385] = ~(t[322] & t[397]);
  assign t[386] = t[398] ^ t[394];
  assign t[387] = ~(t[325] & t[399]);
  assign t[388] = t[400] ^ t[387];
  assign t[389] = t[41] | t[416];
  assign t[38] = ~(t[45] ^ t[63]);
  assign t[390] = t[30] ? x[164] : x[163];
  assign t[391] = ~(t[329] & t[401]);
  assign t[392] = ~(t[331] & t[402]);
  assign t[393] = t[403] ^ t[404];
  assign t[394] = ~(t[335] & t[405]);
  assign t[395] = t[406] ^ t[407];
  assign t[396] = t[57] | t[419];
  assign t[397] = t[61] | t[420];
  assign t[398] = t[413] ? x[166] : x[165];
  assign t[399] = t[64] | t[421];
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[413] ? x[168] : x[167];
  assign t[401] = t[70] | t[424];
  assign t[402] = t[78] | t[426];
  assign t[403] = t[30] ? x[170] : x[169];
  assign t[404] = ~(t[346] & t[408]);
  assign t[405] = t[74] | t[425];
  assign t[406] = t[250] ? x[172] : x[171];
  assign t[407] = ~(t[349] & t[409]);
  assign t[408] = t[123] | t[442];
  assign t[409] = t[116] | t[439];
  assign t[40] = ~(t[39] ^ t[66]);
  assign t[410] = (t[458]);
  assign t[411] = (t[459]);
  assign t[412] = (t[460]);
  assign t[413] = (t[461]);
  assign t[414] = (t[462]);
  assign t[415] = (t[463]);
  assign t[416] = (t[464]);
  assign t[417] = (t[465]);
  assign t[418] = (t[466]);
  assign t[419] = (t[467]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[420] = (t[468]);
  assign t[421] = (t[469]);
  assign t[422] = (t[470]);
  assign t[423] = (t[471]);
  assign t[424] = (t[472]);
  assign t[425] = (t[473]);
  assign t[426] = (t[474]);
  assign t[427] = (t[475]);
  assign t[428] = (t[476]);
  assign t[429] = (t[477]);
  assign t[42] = ~(t[416] | t[69]);
  assign t[430] = (t[478]);
  assign t[431] = (t[479]);
  assign t[432] = (t[480]);
  assign t[433] = (t[481]);
  assign t[434] = (t[482]);
  assign t[435] = (t[483]);
  assign t[436] = (t[484]);
  assign t[437] = (t[485]);
  assign t[438] = (t[486]);
  assign t[439] = (t[487]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (t[488]);
  assign t[441] = (t[489]);
  assign t[442] = (t[490]);
  assign t[443] = (t[491]);
  assign t[444] = (t[492]);
  assign t[445] = (t[493]);
  assign t[446] = (t[494]);
  assign t[447] = (t[495]);
  assign t[448] = (t[496]);
  assign t[449] = (t[497]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (t[498]);
  assign t[451] = (t[499]);
  assign t[452] = (t[500]);
  assign t[453] = (t[501]);
  assign t[454] = (t[502]);
  assign t[455] = (t[503]);
  assign t[456] = (t[504]);
  assign t[457] = (t[505]);
  assign t[458] = t[506] ^ x[5];
  assign t[459] = t[507] ^ x[13];
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = t[508] ^ x[16];
  assign t[461] = t[509] ^ x[19];
  assign t[462] = t[510] ^ x[22];
  assign t[463] = t[511] ^ x[28];
  assign t[464] = t[512] ^ x[34];
  assign t[465] = t[513] ^ x[35];
  assign t[466] = t[514] ^ x[36];
  assign t[467] = t[515] ^ x[42];
  assign t[468] = t[516] ^ x[50];
  assign t[469] = t[517] ^ x[56];
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[470] = t[518] ^ x[57];
  assign t[471] = t[519] ^ x[58];
  assign t[472] = t[520] ^ x[64];
  assign t[473] = t[521] ^ x[72];
  assign t[474] = t[522] ^ x[78];
  assign t[475] = t[523] ^ x[79];
  assign t[476] = t[524] ^ x[80];
  assign t[477] = t[525] ^ x[81];
  assign t[478] = t[526] ^ x[82];
  assign t[479] = t[527] ^ x[83];
  assign t[47] = ~(t[78] | t[79]);
  assign t[480] = t[528] ^ x[86];
  assign t[481] = t[529] ^ x[87];
  assign t[482] = t[530] ^ x[90];
  assign t[483] = t[531] ^ x[91];
  assign t[484] = t[532] ^ x[92];
  assign t[485] = t[533] ^ x[93];
  assign t[486] = t[534] ^ x[94];
  assign t[487] = t[535] ^ x[100];
  assign t[488] = t[536] ^ x[103];
  assign t[489] = t[537] ^ x[104];
  assign t[48] = ~(t[80] ^ t[81]);
  assign t[490] = t[538] ^ x[110];
  assign t[491] = t[539] ^ x[113];
  assign t[492] = t[540] ^ x[114];
  assign t[493] = t[541] ^ x[115];
  assign t[494] = t[542] ^ x[116];
  assign t[495] = t[543] ^ x[117];
  assign t[496] = t[544] ^ x[118];
  assign t[497] = t[545] ^ x[119];
  assign t[498] = t[546] ^ x[120];
  assign t[499] = t[547] ^ x[121];
  assign t[49] = ~(t[413]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = t[548] ^ x[122];
  assign t[501] = t[549] ^ x[123];
  assign t[502] = t[550] ^ x[124];
  assign t[503] = t[551] ^ x[125];
  assign t[504] = t[552] ^ x[141];
  assign t[505] = t[553] ^ x[157];
  assign t[506] = (~t[554] & t[555]);
  assign t[507] = (~t[556] & t[557]);
  assign t[508] = (~t[558] & t[559]);
  assign t[509] = (~t[560] & t[561]);
  assign t[50] = ~(t[82] | t[83]);
  assign t[510] = (~t[562] & t[563]);
  assign t[511] = (~t[564] & t[565]);
  assign t[512] = (~t[566] & t[567]);
  assign t[513] = (~t[564] & t[568]);
  assign t[514] = (~t[564] & t[569]);
  assign t[515] = (~t[570] & t[571]);
  assign t[516] = (~t[572] & t[573]);
  assign t[517] = (~t[574] & t[575]);
  assign t[518] = (~t[566] & t[576]);
  assign t[519] = (~t[566] & t[577]);
  assign t[51] = ~(t[82] | t[84]);
  assign t[520] = (~t[578] & t[579]);
  assign t[521] = (~t[580] & t[581]);
  assign t[522] = (~t[582] & t[583]);
  assign t[523] = (~t[564] & t[584]);
  assign t[524] = (~t[570] & t[585]);
  assign t[525] = (~t[570] & t[586]);
  assign t[526] = (~t[572] & t[587]);
  assign t[527] = (~t[572] & t[588]);
  assign t[528] = (~t[574] & t[589]);
  assign t[529] = (~t[574] & t[590]);
  assign t[52] = t[85] | t[86];
  assign t[530] = (~t[566] & t[591]);
  assign t[531] = (~t[578] & t[592]);
  assign t[532] = (~t[578] & t[593]);
  assign t[533] = (~t[580] & t[594]);
  assign t[534] = (~t[580] & t[595]);
  assign t[535] = (~t[596] & t[597]);
  assign t[536] = (~t[582] & t[598]);
  assign t[537] = (~t[582] & t[599]);
  assign t[538] = (~t[600] & t[601]);
  assign t[539] = (~t[570] & t[602]);
  assign t[53] = ~(t[87] & t[88]);
  assign t[540] = (~t[572] & t[603]);
  assign t[541] = (~t[574] & t[604]);
  assign t[542] = (~t[578] & t[605]);
  assign t[543] = (~t[580] & t[606]);
  assign t[544] = (~t[596] & t[607]);
  assign t[545] = (~t[596] & t[608]);
  assign t[546] = (~t[582] & t[609]);
  assign t[547] = (~t[600] & t[610]);
  assign t[548] = (~t[600] & t[611]);
  assign t[549] = (~t[596] & t[612]);
  assign t[54] = ~(t[417]);
  assign t[550] = (~t[600] & t[613]);
  assign t[551] = (~t[554] & t[614]);
  assign t[552] = (~t[554] & t[615]);
  assign t[553] = (~t[554] & t[616]);
  assign t[554] = t[617] ^ x[4];
  assign t[555] = t[618] ^ x[5];
  assign t[556] = t[619] ^ x[12];
  assign t[557] = t[620] ^ x[13];
  assign t[558] = t[621] ^ x[15];
  assign t[559] = t[622] ^ x[16];
  assign t[55] = ~(t[418]);
  assign t[560] = t[623] ^ x[18];
  assign t[561] = t[624] ^ x[19];
  assign t[562] = t[625] ^ x[21];
  assign t[563] = t[626] ^ x[22];
  assign t[564] = t[627] ^ x[27];
  assign t[565] = t[628] ^ x[28];
  assign t[566] = t[629] ^ x[33];
  assign t[567] = t[630] ^ x[34];
  assign t[568] = t[631] ^ x[35];
  assign t[569] = t[632] ^ x[36];
  assign t[56] = ~(t[89] | t[90]);
  assign t[570] = t[633] ^ x[41];
  assign t[571] = t[634] ^ x[42];
  assign t[572] = t[635] ^ x[49];
  assign t[573] = t[636] ^ x[50];
  assign t[574] = t[637] ^ x[55];
  assign t[575] = t[638] ^ x[56];
  assign t[576] = t[639] ^ x[57];
  assign t[577] = t[640] ^ x[58];
  assign t[578] = t[641] ^ x[63];
  assign t[579] = t[642] ^ x[64];
  assign t[57] = ~(t[91] | t[92]);
  assign t[580] = t[643] ^ x[71];
  assign t[581] = t[644] ^ x[72];
  assign t[582] = t[645] ^ x[77];
  assign t[583] = t[646] ^ x[78];
  assign t[584] = t[647] ^ x[79];
  assign t[585] = t[648] ^ x[80];
  assign t[586] = t[649] ^ x[81];
  assign t[587] = t[650] ^ x[82];
  assign t[588] = t[651] ^ x[83];
  assign t[589] = t[652] ^ x[86];
  assign t[58] = ~(t[419] | t[93]);
  assign t[590] = t[653] ^ x[87];
  assign t[591] = t[654] ^ x[90];
  assign t[592] = t[655] ^ x[91];
  assign t[593] = t[656] ^ x[92];
  assign t[594] = t[657] ^ x[93];
  assign t[595] = t[658] ^ x[94];
  assign t[596] = t[659] ^ x[99];
  assign t[597] = t[660] ^ x[100];
  assign t[598] = t[661] ^ x[103];
  assign t[599] = t[662] ^ x[104];
  assign t[59] = t[413] ? x[44] : x[43];
  assign t[5] = t[9] ^ x[8];
  assign t[600] = t[663] ^ x[109];
  assign t[601] = t[664] ^ x[110];
  assign t[602] = t[665] ^ x[113];
  assign t[603] = t[666] ^ x[114];
  assign t[604] = t[667] ^ x[115];
  assign t[605] = t[668] ^ x[116];
  assign t[606] = t[669] ^ x[117];
  assign t[607] = t[670] ^ x[118];
  assign t[608] = t[671] ^ x[119];
  assign t[609] = t[672] ^ x[120];
  assign t[60] = ~(t[94] & t[95]);
  assign t[610] = t[673] ^ x[121];
  assign t[611] = t[674] ^ x[122];
  assign t[612] = t[675] ^ x[123];
  assign t[613] = t[676] ^ x[124];
  assign t[614] = t[677] ^ x[125];
  assign t[615] = t[678] ^ x[141];
  assign t[616] = t[679] ^ x[157];
  assign t[617] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[618] = (x[0]);
  assign t[619] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = ~(t[96] | t[97]);
  assign t[620] = (x[11]);
  assign t[621] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[622] = (x[14]);
  assign t[623] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[624] = (x[17]);
  assign t[625] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[626] = (x[20]);
  assign t[627] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[628] = (x[24]);
  assign t[629] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[62] = ~(t[420] | t[98]);
  assign t[630] = (x[30]);
  assign t[631] = (x[25]);
  assign t[632] = (x[26]);
  assign t[633] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[634] = (x[38]);
  assign t[635] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[636] = (x[46]);
  assign t[637] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[638] = (x[52]);
  assign t[639] = (x[31]);
  assign t[63] = ~(t[99] ^ t[100]);
  assign t[640] = (x[32]);
  assign t[641] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[642] = (x[60]);
  assign t[643] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[644] = (x[68]);
  assign t[645] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[646] = (x[74]);
  assign t[647] = (x[23]);
  assign t[648] = (x[39]);
  assign t[649] = (x[40]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[650] = (x[47]);
  assign t[651] = (x[48]);
  assign t[652] = (x[53]);
  assign t[653] = (x[54]);
  assign t[654] = (x[29]);
  assign t[655] = (x[61]);
  assign t[656] = (x[62]);
  assign t[657] = (x[69]);
  assign t[658] = (x[70]);
  assign t[659] = (x[95] & ~x[96] & ~x[97] & ~x[98]) | (~x[95] & x[96] & ~x[97] & ~x[98]) | (~x[95] & ~x[96] & x[97] & ~x[98]) | (~x[95] & ~x[96] & ~x[97] & x[98]) | (x[95] & x[96] & x[97] & ~x[98]) | (x[95] & x[96] & ~x[97] & x[98]) | (x[95] & ~x[96] & x[97] & x[98]) | (~x[95] & x[96] & x[97] & x[98]);
  assign t[65] = ~(t[421] | t[103]);
  assign t[660] = (x[96]);
  assign t[661] = (x[75]);
  assign t[662] = (x[76]);
  assign t[663] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[664] = (x[106]);
  assign t[665] = (x[37]);
  assign t[666] = (x[45]);
  assign t[667] = (x[51]);
  assign t[668] = (x[59]);
  assign t[669] = (x[67]);
  assign t[66] = ~(t[104] ^ t[105]);
  assign t[670] = (x[97]);
  assign t[671] = (x[98]);
  assign t[672] = (x[73]);
  assign t[673] = (x[107]);
  assign t[674] = (x[108]);
  assign t[675] = (x[95]);
  assign t[676] = (x[105]);
  assign t[677] = (x[1]);
  assign t[678] = (x[2]);
  assign t[679] = (x[3]);
  assign t[67] = ~(t[422]);
  assign t[68] = ~(t[423]);
  assign t[69] = ~(t[106] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[424] | t[110]);
  assign t[72] = t[30] ? x[66] : x[65];
  assign t[73] = ~(t[111] & t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[425] | t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[120] | t[121]);
  assign t[79] = ~(t[426] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[123] | t[124]);
  assign t[81] = ~(t[125] ^ t[126]);
  assign t[82] = ~(t[127]);
  assign t[83] = t[411] ? t[129] : t[128];
  assign t[84] = t[411] ? t[131] : t[130];
  assign t[85] = ~(t[132] & t[133]);
  assign t[86] = ~(t[82] | t[134]);
  assign t[87] = ~(t[135] | t[136]);
  assign t[88] = t[127] | t[137];
  assign t[89] = ~(t[427]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[417] | t[418]);
  assign t[91] = ~(t[428]);
  assign t[92] = ~(t[429]);
  assign t[93] = ~(t[138] | t[139]);
  assign t[94] = ~(t[140] | t[141]);
  assign t[95] = ~(t[142] | t[143]);
  assign t[96] = ~(t[430]);
  assign t[97] = ~(t[431]);
  assign t[98] = ~(t[144] | t[145]);
  assign t[99] = t[146] ? x[85] : x[84];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[212] & ~t[282] & ~t[361]) | (~t[0] & t[212] & ~t[282] & ~t[361]) | (~t[0] & ~t[212] & t[282] & ~t[361]) | (~t[0] & ~t[212] & ~t[282] & t[361]) | (t[0] & t[212] & t[282] & ~t[361]) | (t[0] & t[212] & ~t[282] & t[361]) | (t[0] & ~t[212] & t[282] & t[361]) | (~t[0] & t[212] & t[282] & t[361]);
endmodule

module R2ind146(x, y);
 input [124:0] x;
 output y;

 wire [364:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[149]);
  assign t[103] = ~(t[108] | t[101]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[5];
  assign t[156] = t[201] ^ x[13];
  assign t[157] = t[202] ^ x[16];
  assign t[158] = t[203] ^ x[19];
  assign t[159] = t[204] ^ x[22];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[28];
  assign t[161] = t[206] ^ x[36];
  assign t[162] = t[207] ^ x[39];
  assign t[163] = t[208] ^ x[40];
  assign t[164] = t[209] ^ x[46];
  assign t[165] = t[210] ^ x[52];
  assign t[166] = t[211] ^ x[60];
  assign t[167] = t[212] ^ x[63];
  assign t[168] = t[213] ^ x[64];
  assign t[169] = t[214] ^ x[70];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[76];
  assign t[171] = t[216] ^ x[84];
  assign t[172] = t[217] ^ x[87];
  assign t[173] = t[218] ^ x[88];
  assign t[174] = t[219] ^ x[89];
  assign t[175] = t[220] ^ x[90];
  assign t[176] = t[221] ^ x[91];
  assign t[177] = t[222] ^ x[92];
  assign t[178] = t[223] ^ x[93];
  assign t[179] = t[224] ^ x[94];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[95];
  assign t[181] = t[226] ^ x[96];
  assign t[182] = t[227] ^ x[97];
  assign t[183] = t[228] ^ x[98];
  assign t[184] = t[229] ^ x[104];
  assign t[185] = t[230] ^ x[105];
  assign t[186] = t[231] ^ x[106];
  assign t[187] = t[232] ^ x[112];
  assign t[188] = t[233] ^ x[113];
  assign t[189] = t[234] ^ x[114];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[115];
  assign t[191] = t[236] ^ x[116];
  assign t[192] = t[237] ^ x[117];
  assign t[193] = t[238] ^ x[118];
  assign t[194] = t[239] ^ x[119];
  assign t[195] = t[240] ^ x[120];
  assign t[196] = t[241] ^ x[121];
  assign t[197] = t[242] ^ x[122];
  assign t[198] = t[243] ^ x[123];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[245] & t[246]);
  assign t[201] = (~t[247] & t[248]);
  assign t[202] = (~t[249] & t[250]);
  assign t[203] = (~t[251] & t[252]);
  assign t[204] = (~t[253] & t[254]);
  assign t[205] = (~t[255] & t[256]);
  assign t[206] = (~t[257] & t[258]);
  assign t[207] = (~t[255] & t[259]);
  assign t[208] = (~t[255] & t[260]);
  assign t[209] = (~t[261] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[263] & t[264]);
  assign t[211] = (~t[265] & t[266]);
  assign t[212] = (~t[257] & t[267]);
  assign t[213] = (~t[257] & t[268]);
  assign t[214] = (~t[269] & t[270]);
  assign t[215] = (~t[271] & t[272]);
  assign t[216] = (~t[273] & t[274]);
  assign t[217] = (~t[255] & t[275]);
  assign t[218] = (~t[261] & t[276]);
  assign t[219] = (~t[261] & t[277]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[263] & t[278]);
  assign t[221] = (~t[263] & t[279]);
  assign t[222] = (~t[265] & t[280]);
  assign t[223] = (~t[265] & t[281]);
  assign t[224] = (~t[257] & t[282]);
  assign t[225] = (~t[269] & t[283]);
  assign t[226] = (~t[269] & t[284]);
  assign t[227] = (~t[271] & t[285]);
  assign t[228] = (~t[271] & t[286]);
  assign t[229] = (~t[287] & t[288]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[273] & t[289]);
  assign t[231] = (~t[273] & t[290]);
  assign t[232] = (~t[291] & t[292]);
  assign t[233] = (~t[261] & t[293]);
  assign t[234] = (~t[263] & t[294]);
  assign t[235] = (~t[265] & t[295]);
  assign t[236] = (~t[269] & t[296]);
  assign t[237] = (~t[271] & t[297]);
  assign t[238] = (~t[287] & t[298]);
  assign t[239] = (~t[287] & t[299]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[273] & t[300]);
  assign t[241] = (~t[291] & t[301]);
  assign t[242] = (~t[291] & t[302]);
  assign t[243] = (~t[287] & t[303]);
  assign t[244] = (~t[291] & t[304]);
  assign t[245] = t[305] ^ x[4];
  assign t[246] = t[306] ^ x[5];
  assign t[247] = t[307] ^ x[12];
  assign t[248] = t[308] ^ x[13];
  assign t[249] = t[309] ^ x[15];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[310] ^ x[16];
  assign t[251] = t[311] ^ x[18];
  assign t[252] = t[312] ^ x[19];
  assign t[253] = t[313] ^ x[21];
  assign t[254] = t[314] ^ x[22];
  assign t[255] = t[315] ^ x[27];
  assign t[256] = t[316] ^ x[28];
  assign t[257] = t[317] ^ x[35];
  assign t[258] = t[318] ^ x[36];
  assign t[259] = t[319] ^ x[39];
  assign t[25] = ~(t[113]);
  assign t[260] = t[320] ^ x[40];
  assign t[261] = t[321] ^ x[45];
  assign t[262] = t[322] ^ x[46];
  assign t[263] = t[323] ^ x[51];
  assign t[264] = t[324] ^ x[52];
  assign t[265] = t[325] ^ x[59];
  assign t[266] = t[326] ^ x[60];
  assign t[267] = t[327] ^ x[63];
  assign t[268] = t[328] ^ x[64];
  assign t[269] = t[329] ^ x[69];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[70];
  assign t[271] = t[331] ^ x[75];
  assign t[272] = t[332] ^ x[76];
  assign t[273] = t[333] ^ x[83];
  assign t[274] = t[334] ^ x[84];
  assign t[275] = t[335] ^ x[87];
  assign t[276] = t[336] ^ x[88];
  assign t[277] = t[337] ^ x[89];
  assign t[278] = t[338] ^ x[90];
  assign t[279] = t[339] ^ x[91];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[92];
  assign t[281] = t[341] ^ x[93];
  assign t[282] = t[342] ^ x[94];
  assign t[283] = t[343] ^ x[95];
  assign t[284] = t[344] ^ x[96];
  assign t[285] = t[345] ^ x[97];
  assign t[286] = t[346] ^ x[98];
  assign t[287] = t[347] ^ x[103];
  assign t[288] = t[348] ^ x[104];
  assign t[289] = t[349] ^ x[105];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[106];
  assign t[291] = t[351] ^ x[111];
  assign t[292] = t[352] ^ x[112];
  assign t[293] = t[353] ^ x[113];
  assign t[294] = t[354] ^ x[114];
  assign t[295] = t[355] ^ x[115];
  assign t[296] = t[356] ^ x[116];
  assign t[297] = t[357] ^ x[117];
  assign t[298] = t[358] ^ x[118];
  assign t[299] = t[359] ^ x[119];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[120];
  assign t[301] = t[361] ^ x[121];
  assign t[302] = t[362] ^ x[122];
  assign t[303] = t[363] ^ x[123];
  assign t[304] = t[364] ^ x[124];
  assign t[305] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[306] = (x[3]);
  assign t[307] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[308] = (x[11]);
  assign t[309] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = (x[14]);
  assign t[311] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[312] = (x[17]);
  assign t[313] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[314] = (x[20]);
  assign t[315] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[316] = (x[24]);
  assign t[317] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[318] = (x[32]);
  assign t[319] = (x[26]);
  assign t[31] = t[48] | t[115];
  assign t[320] = (x[23]);
  assign t[321] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[322] = (x[42]);
  assign t[323] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[324] = (x[48]);
  assign t[325] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[326] = (x[56]);
  assign t[327] = (x[34]);
  assign t[328] = (x[31]);
  assign t[329] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[32] = t[49] ? x[30] : x[29];
  assign t[330] = (x[66]);
  assign t[331] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[332] = (x[72]);
  assign t[333] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[334] = (x[80]);
  assign t[335] = (x[25]);
  assign t[336] = (x[44]);
  assign t[337] = (x[41]);
  assign t[338] = (x[50]);
  assign t[339] = (x[47]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[58]);
  assign t[341] = (x[55]);
  assign t[342] = (x[33]);
  assign t[343] = (x[68]);
  assign t[344] = (x[65]);
  assign t[345] = (x[74]);
  assign t[346] = (x[71]);
  assign t[347] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[348] = (x[100]);
  assign t[349] = (x[82]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[79]);
  assign t[351] = (x[107] & ~x[108] & ~x[109] & ~x[110]) | (~x[107] & x[108] & ~x[109] & ~x[110]) | (~x[107] & ~x[108] & x[109] & ~x[110]) | (~x[107] & ~x[108] & ~x[109] & x[110]) | (x[107] & x[108] & x[109] & ~x[110]) | (x[107] & x[108] & ~x[109] & x[110]) | (x[107] & ~x[108] & x[109] & x[110]) | (~x[107] & x[108] & x[109] & x[110]);
  assign t[352] = (x[108]);
  assign t[353] = (x[43]);
  assign t[354] = (x[49]);
  assign t[355] = (x[57]);
  assign t[356] = (x[67]);
  assign t[357] = (x[73]);
  assign t[358] = (x[102]);
  assign t[359] = (x[99]);
  assign t[35] = t[54] ^ t[44];
  assign t[360] = (x[81]);
  assign t[361] = (x[110]);
  assign t[362] = (x[107]);
  assign t[363] = (x[101]);
  assign t[364] = (x[109]);
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[36];
  assign t[38] = ~(t[58] & t[59]);
  assign t[39] = t[60] | t[116];
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[38] : x[37];
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[119];
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = t[77] | t[120];
  assign t[54] = t[113] ? x[54] : x[53];
  assign t[55] = ~(t[78] & t[79]);
  assign t[56] = t[80] | t[121];
  assign t[57] = t[113] ? x[62] : x[61];
  assign t[58] = ~(t[122]);
  assign t[59] = ~(t[123]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[81] | t[58]);
  assign t[61] = ~(t[82] & t[83]);
  assign t[62] = t[84] | t[124];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = t[87] | t[125];
  assign t[65] = t[18] ? x[78] : x[77];
  assign t[66] = ~(t[88] & t[89]);
  assign t[67] = ~(t[90] & t[91]);
  assign t[68] = t[92] | t[126];
  assign t[69] = t[93] ? x[86] : x[85];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[94] & t[95]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[98] | t[78]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[101] & t[102]);
  assign t[89] = t[103] | t[139];
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[140]);
  assign t[91] = ~(t[141]);
  assign t[92] = ~(t[104] | t[90]);
  assign t[93] = ~(t[25]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [124:0] x;
 output y;

 wire [373:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[142] & t[141]);
  assign t[102] = ~(t[154]);
  assign t[103] = ~(t[145] & t[144]);
  assign t[104] = ~(t[155]);
  assign t[105] = ~(t[147] & t[146]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[158]);
  assign t[109] = ~(t[115] & t[116]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[117] & t[118]);
  assign t[115] = ~(t[158] & t[157]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[161] & t[160]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[5];
  assign t[165] = t[210] ^ x[13];
  assign t[166] = t[211] ^ x[16];
  assign t[167] = t[212] ^ x[19];
  assign t[168] = t[213] ^ x[22];
  assign t[169] = t[214] ^ x[28];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[36];
  assign t[171] = t[216] ^ x[39];
  assign t[172] = t[217] ^ x[40];
  assign t[173] = t[218] ^ x[46];
  assign t[174] = t[219] ^ x[52];
  assign t[175] = t[220] ^ x[60];
  assign t[176] = t[221] ^ x[63];
  assign t[177] = t[222] ^ x[64];
  assign t[178] = t[223] ^ x[70];
  assign t[179] = t[224] ^ x[76];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[84];
  assign t[181] = t[226] ^ x[87];
  assign t[182] = t[227] ^ x[88];
  assign t[183] = t[228] ^ x[89];
  assign t[184] = t[229] ^ x[90];
  assign t[185] = t[230] ^ x[91];
  assign t[186] = t[231] ^ x[92];
  assign t[187] = t[232] ^ x[93];
  assign t[188] = t[233] ^ x[94];
  assign t[189] = t[234] ^ x[95];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[96];
  assign t[191] = t[236] ^ x[97];
  assign t[192] = t[237] ^ x[98];
  assign t[193] = t[238] ^ x[104];
  assign t[194] = t[239] ^ x[105];
  assign t[195] = t[240] ^ x[106];
  assign t[196] = t[241] ^ x[112];
  assign t[197] = t[242] ^ x[113];
  assign t[198] = t[243] ^ x[114];
  assign t[199] = t[244] ^ x[115];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[116];
  assign t[201] = t[246] ^ x[117];
  assign t[202] = t[247] ^ x[118];
  assign t[203] = t[248] ^ x[119];
  assign t[204] = t[249] ^ x[120];
  assign t[205] = t[250] ^ x[121];
  assign t[206] = t[251] ^ x[122];
  assign t[207] = t[252] ^ x[123];
  assign t[208] = t[253] ^ x[124];
  assign t[209] = (~t[254] & t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[256] & t[257]);
  assign t[211] = (~t[258] & t[259]);
  assign t[212] = (~t[260] & t[261]);
  assign t[213] = (~t[262] & t[263]);
  assign t[214] = (~t[264] & t[265]);
  assign t[215] = (~t[266] & t[267]);
  assign t[216] = (~t[264] & t[268]);
  assign t[217] = (~t[264] & t[269]);
  assign t[218] = (~t[270] & t[271]);
  assign t[219] = (~t[272] & t[273]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[274] & t[275]);
  assign t[221] = (~t[266] & t[276]);
  assign t[222] = (~t[266] & t[277]);
  assign t[223] = (~t[278] & t[279]);
  assign t[224] = (~t[280] & t[281]);
  assign t[225] = (~t[282] & t[283]);
  assign t[226] = (~t[264] & t[284]);
  assign t[227] = (~t[270] & t[285]);
  assign t[228] = (~t[270] & t[286]);
  assign t[229] = (~t[272] & t[287]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[272] & t[288]);
  assign t[231] = (~t[274] & t[289]);
  assign t[232] = (~t[274] & t[290]);
  assign t[233] = (~t[266] & t[291]);
  assign t[234] = (~t[278] & t[292]);
  assign t[235] = (~t[278] & t[293]);
  assign t[236] = (~t[280] & t[294]);
  assign t[237] = (~t[280] & t[295]);
  assign t[238] = (~t[296] & t[297]);
  assign t[239] = (~t[282] & t[298]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[282] & t[299]);
  assign t[241] = (~t[300] & t[301]);
  assign t[242] = (~t[270] & t[302]);
  assign t[243] = (~t[272] & t[303]);
  assign t[244] = (~t[274] & t[304]);
  assign t[245] = (~t[278] & t[305]);
  assign t[246] = (~t[280] & t[306]);
  assign t[247] = (~t[296] & t[307]);
  assign t[248] = (~t[296] & t[308]);
  assign t[249] = (~t[282] & t[309]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = (~t[300] & t[310]);
  assign t[251] = (~t[300] & t[311]);
  assign t[252] = (~t[296] & t[312]);
  assign t[253] = (~t[300] & t[313]);
  assign t[254] = t[314] ^ x[4];
  assign t[255] = t[315] ^ x[5];
  assign t[256] = t[316] ^ x[12];
  assign t[257] = t[317] ^ x[13];
  assign t[258] = t[318] ^ x[15];
  assign t[259] = t[319] ^ x[16];
  assign t[25] = ~(t[122]);
  assign t[260] = t[320] ^ x[18];
  assign t[261] = t[321] ^ x[19];
  assign t[262] = t[322] ^ x[21];
  assign t[263] = t[323] ^ x[22];
  assign t[264] = t[324] ^ x[27];
  assign t[265] = t[325] ^ x[28];
  assign t[266] = t[326] ^ x[35];
  assign t[267] = t[327] ^ x[36];
  assign t[268] = t[328] ^ x[39];
  assign t[269] = t[329] ^ x[40];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[45];
  assign t[271] = t[331] ^ x[46];
  assign t[272] = t[332] ^ x[51];
  assign t[273] = t[333] ^ x[52];
  assign t[274] = t[334] ^ x[59];
  assign t[275] = t[335] ^ x[60];
  assign t[276] = t[336] ^ x[63];
  assign t[277] = t[337] ^ x[64];
  assign t[278] = t[338] ^ x[69];
  assign t[279] = t[339] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[75];
  assign t[281] = t[341] ^ x[76];
  assign t[282] = t[342] ^ x[83];
  assign t[283] = t[343] ^ x[84];
  assign t[284] = t[344] ^ x[87];
  assign t[285] = t[345] ^ x[88];
  assign t[286] = t[346] ^ x[89];
  assign t[287] = t[347] ^ x[90];
  assign t[288] = t[348] ^ x[91];
  assign t[289] = t[349] ^ x[92];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[93];
  assign t[291] = t[351] ^ x[94];
  assign t[292] = t[352] ^ x[95];
  assign t[293] = t[353] ^ x[96];
  assign t[294] = t[354] ^ x[97];
  assign t[295] = t[355] ^ x[98];
  assign t[296] = t[356] ^ x[103];
  assign t[297] = t[357] ^ x[104];
  assign t[298] = t[358] ^ x[105];
  assign t[299] = t[359] ^ x[106];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[111];
  assign t[301] = t[361] ^ x[112];
  assign t[302] = t[362] ^ x[113];
  assign t[303] = t[363] ^ x[114];
  assign t[304] = t[364] ^ x[115];
  assign t[305] = t[365] ^ x[116];
  assign t[306] = t[366] ^ x[117];
  assign t[307] = t[367] ^ x[118];
  assign t[308] = t[368] ^ x[119];
  assign t[309] = t[369] ^ x[120];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[370] ^ x[121];
  assign t[311] = t[371] ^ x[122];
  assign t[312] = t[372] ^ x[123];
  assign t[313] = t[373] ^ x[124];
  assign t[314] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[315] = (x[2]);
  assign t[316] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[317] = (x[11]);
  assign t[318] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[319] = (x[14]);
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[321] = (x[17]);
  assign t[322] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[323] = (x[20]);
  assign t[324] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[325] = (x[24]);
  assign t[326] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[327] = (x[32]);
  assign t[328] = (x[26]);
  assign t[329] = (x[23]);
  assign t[32] = t[18] ? x[30] : x[29];
  assign t[330] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[331] = (x[42]);
  assign t[332] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[333] = (x[48]);
  assign t[334] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[335] = (x[56]);
  assign t[336] = (x[34]);
  assign t[337] = (x[31]);
  assign t[338] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[339] = (x[66]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[341] = (x[72]);
  assign t[342] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[343] = (x[80]);
  assign t[344] = (x[25]);
  assign t[345] = (x[44]);
  assign t[346] = (x[41]);
  assign t[347] = (x[50]);
  assign t[348] = (x[47]);
  assign t[349] = (x[58]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[55]);
  assign t[351] = (x[33]);
  assign t[352] = (x[68]);
  assign t[353] = (x[65]);
  assign t[354] = (x[74]);
  assign t[355] = (x[71]);
  assign t[356] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[357] = (x[100]);
  assign t[358] = (x[82]);
  assign t[359] = (x[79]);
  assign t[35] = t[53] ^ t[44];
  assign t[360] = (x[107] & ~x[108] & ~x[109] & ~x[110]) | (~x[107] & x[108] & ~x[109] & ~x[110]) | (~x[107] & ~x[108] & x[109] & ~x[110]) | (~x[107] & ~x[108] & ~x[109] & x[110]) | (x[107] & x[108] & x[109] & ~x[110]) | (x[107] & x[108] & ~x[109] & x[110]) | (x[107] & ~x[108] & x[109] & x[110]) | (~x[107] & x[108] & x[109] & x[110]);
  assign t[361] = (x[108]);
  assign t[362] = (x[43]);
  assign t[363] = (x[49]);
  assign t[364] = (x[57]);
  assign t[365] = (x[67]);
  assign t[366] = (x[73]);
  assign t[367] = (x[102]);
  assign t[368] = (x[99]);
  assign t[369] = (x[81]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[370] = (x[110]);
  assign t[371] = (x[107]);
  assign t[372] = (x[101]);
  assign t[373] = (x[109]);
  assign t[37] = t[56] ^ t[36];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = ~(t[59] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[122] ? x[38] : x[37];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = ~(t[72] & t[73]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[74] & t[128]);
  assign t[51] = ~(t[75] & t[76]);
  assign t[52] = ~(t[77] & t[129]);
  assign t[53] = t[122] ? x[54] : x[53];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = ~(t[80] & t[130]);
  assign t[56] = t[122] ? x[62] : x[61];
  assign t[57] = ~(t[131]);
  assign t[58] = ~(t[132]);
  assign t[59] = ~(t[81] & t[82]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[83] & t[84]);
  assign t[61] = ~(t[85] & t[133]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[134]);
  assign t[64] = t[18] ? x[78] : x[77];
  assign t[65] = ~(t[89] & t[90]);
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = ~(t[93] & t[135]);
  assign t[68] = t[94] ? x[86] : x[85];
  assign t[69] = ~(t[95] & t[96]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[127] & t[126]);
  assign t[71] = ~(t[136]);
  assign t[72] = ~(t[137]);
  assign t[73] = ~(t[138]);
  assign t[74] = ~(t[97] & t[98]);
  assign t[75] = ~(t[139]);
  assign t[76] = ~(t[140]);
  assign t[77] = ~(t[99] & t[100]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[142]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[101] & t[102]);
  assign t[81] = ~(t[132] & t[131]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[145]);
  assign t[85] = ~(t[103] & t[104]);
  assign t[86] = ~(t[146]);
  assign t[87] = ~(t[147]);
  assign t[88] = ~(t[105] & t[106]);
  assign t[89] = ~(t[107] & t[108]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[109] & t[148]);
  assign t[91] = ~(t[149]);
  assign t[92] = ~(t[150]);
  assign t[93] = ~(t[110] & t[111]);
  assign t[94] = ~(t[25]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[114] & t[151]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [114:0] x;
 output y;

 wire [304:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[5];
  assign t[136] = t[171] ^ x[13];
  assign t[137] = t[172] ^ x[16];
  assign t[138] = t[173] ^ x[19];
  assign t[139] = t[174] ^ x[22];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[28];
  assign t[141] = t[176] ^ x[29];
  assign t[142] = t[177] ^ x[37];
  assign t[143] = t[178] ^ x[38];
  assign t[144] = t[179] ^ x[41];
  assign t[145] = t[180] ^ x[47];
  assign t[146] = t[181] ^ x[48];
  assign t[147] = t[182] ^ x[54];
  assign t[148] = t[183] ^ x[55];
  assign t[149] = t[184] ^ x[63];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[64];
  assign t[151] = t[186] ^ x[67];
  assign t[152] = t[187] ^ x[73];
  assign t[153] = t[188] ^ x[74];
  assign t[154] = t[189] ^ x[80];
  assign t[155] = t[190] ^ x[81];
  assign t[156] = t[191] ^ x[89];
  assign t[157] = t[192] ^ x[90];
  assign t[158] = t[193] ^ x[93];
  assign t[159] = t[194] ^ x[94];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[95];
  assign t[161] = t[196] ^ x[96];
  assign t[162] = t[197] ^ x[97];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[104];
  assign t[165] = t[200] ^ x[105];
  assign t[166] = t[201] ^ x[111];
  assign t[167] = t[202] ^ x[112];
  assign t[168] = t[203] ^ x[113];
  assign t[169] = t[204] ^ x[114];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (~t[205] & t[206]);
  assign t[171] = (~t[207] & t[208]);
  assign t[172] = (~t[209] & t[210]);
  assign t[173] = (~t[211] & t[212]);
  assign t[174] = (~t[213] & t[214]);
  assign t[175] = (~t[215] & t[216]);
  assign t[176] = (~t[215] & t[217]);
  assign t[177] = (~t[218] & t[219]);
  assign t[178] = (~t[218] & t[220]);
  assign t[179] = (~t[215] & t[221]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (~t[222] & t[223]);
  assign t[181] = (~t[222] & t[224]);
  assign t[182] = (~t[225] & t[226]);
  assign t[183] = (~t[225] & t[227]);
  assign t[184] = (~t[228] & t[229]);
  assign t[185] = (~t[228] & t[230]);
  assign t[186] = (~t[218] & t[231]);
  assign t[187] = (~t[232] & t[233]);
  assign t[188] = (~t[232] & t[234]);
  assign t[189] = (~t[235] & t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (~t[235] & t[237]);
  assign t[191] = (~t[238] & t[239]);
  assign t[192] = (~t[238] & t[240]);
  assign t[193] = (~t[222] & t[241]);
  assign t[194] = (~t[225] & t[242]);
  assign t[195] = (~t[228] & t[243]);
  assign t[196] = (~t[232] & t[244]);
  assign t[197] = (~t[235] & t[245]);
  assign t[198] = (~t[246] & t[247]);
  assign t[199] = (~t[246] & t[248]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[238] & t[249]);
  assign t[201] = (~t[250] & t[251]);
  assign t[202] = (~t[250] & t[252]);
  assign t[203] = (~t[246] & t[253]);
  assign t[204] = (~t[250] & t[254]);
  assign t[205] = t[255] ^ x[4];
  assign t[206] = t[256] ^ x[5];
  assign t[207] = t[257] ^ x[12];
  assign t[208] = t[258] ^ x[13];
  assign t[209] = t[259] ^ x[15];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[260] ^ x[16];
  assign t[211] = t[261] ^ x[18];
  assign t[212] = t[262] ^ x[19];
  assign t[213] = t[263] ^ x[21];
  assign t[214] = t[264] ^ x[22];
  assign t[215] = t[265] ^ x[27];
  assign t[216] = t[266] ^ x[28];
  assign t[217] = t[267] ^ x[29];
  assign t[218] = t[268] ^ x[36];
  assign t[219] = t[269] ^ x[37];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[270] ^ x[38];
  assign t[221] = t[271] ^ x[41];
  assign t[222] = t[272] ^ x[46];
  assign t[223] = t[273] ^ x[47];
  assign t[224] = t[274] ^ x[48];
  assign t[225] = t[275] ^ x[53];
  assign t[226] = t[276] ^ x[54];
  assign t[227] = t[277] ^ x[55];
  assign t[228] = t[278] ^ x[62];
  assign t[229] = t[279] ^ x[63];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[280] ^ x[64];
  assign t[231] = t[281] ^ x[67];
  assign t[232] = t[282] ^ x[72];
  assign t[233] = t[283] ^ x[73];
  assign t[234] = t[284] ^ x[74];
  assign t[235] = t[285] ^ x[79];
  assign t[236] = t[286] ^ x[80];
  assign t[237] = t[287] ^ x[81];
  assign t[238] = t[288] ^ x[88];
  assign t[239] = t[289] ^ x[89];
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = t[290] ^ x[90];
  assign t[241] = t[291] ^ x[93];
  assign t[242] = t[292] ^ x[94];
  assign t[243] = t[293] ^ x[95];
  assign t[244] = t[294] ^ x[96];
  assign t[245] = t[295] ^ x[97];
  assign t[246] = t[296] ^ x[102];
  assign t[247] = t[297] ^ x[103];
  assign t[248] = t[298] ^ x[104];
  assign t[249] = t[299] ^ x[105];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[300] ^ x[110];
  assign t[251] = t[301] ^ x[111];
  assign t[252] = t[302] ^ x[112];
  assign t[253] = t[303] ^ x[113];
  assign t[254] = t[304] ^ x[114];
  assign t[255] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[256] = (x[1]);
  assign t[257] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[258] = (x[11]);
  assign t[259] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[25] = ~(t[103]);
  assign t[260] = (x[14]);
  assign t[261] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[262] = (x[17]);
  assign t[263] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[264] = (x[20]);
  assign t[265] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[266] = (x[25]);
  assign t[267] = (x[23]);
  assign t[268] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[269] = (x[34]);
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = (x[32]);
  assign t[271] = (x[26]);
  assign t[272] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[273] = (x[44]);
  assign t[274] = (x[42]);
  assign t[275] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[276] = (x[51]);
  assign t[277] = (x[49]);
  assign t[278] = (x[58] & ~x[59] & ~x[60] & ~x[61]) | (~x[58] & x[59] & ~x[60] & ~x[61]) | (~x[58] & ~x[59] & x[60] & ~x[61]) | (~x[58] & ~x[59] & ~x[60] & x[61]) | (x[58] & x[59] & x[60] & ~x[61]) | (x[58] & x[59] & ~x[60] & x[61]) | (x[58] & ~x[59] & x[60] & x[61]) | (~x[58] & x[59] & x[60] & x[61]);
  assign t[279] = (x[60]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[58]);
  assign t[281] = (x[35]);
  assign t[282] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[283] = (x[70]);
  assign t[284] = (x[68]);
  assign t[285] = (x[75] & ~x[76] & ~x[77] & ~x[78]) | (~x[75] & x[76] & ~x[77] & ~x[78]) | (~x[75] & ~x[76] & x[77] & ~x[78]) | (~x[75] & ~x[76] & ~x[77] & x[78]) | (x[75] & x[76] & x[77] & ~x[78]) | (x[75] & x[76] & ~x[77] & x[78]) | (x[75] & ~x[76] & x[77] & x[78]) | (~x[75] & x[76] & x[77] & x[78]);
  assign t[286] = (x[77]);
  assign t[287] = (x[75]);
  assign t[288] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[289] = (x[86]);
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = (x[84]);
  assign t[291] = (x[45]);
  assign t[292] = (x[52]);
  assign t[293] = (x[61]);
  assign t[294] = (x[71]);
  assign t[295] = (x[78]);
  assign t[296] = (x[98] & ~x[99] & ~x[100] & ~x[101]) | (~x[98] & x[99] & ~x[100] & ~x[101]) | (~x[98] & ~x[99] & x[100] & ~x[101]) | (~x[98] & ~x[99] & ~x[100] & x[101]) | (x[98] & x[99] & x[100] & ~x[101]) | (x[98] & x[99] & ~x[100] & x[101]) | (x[98] & ~x[99] & x[100] & x[101]) | (~x[98] & x[99] & x[100] & x[101]);
  assign t[297] = (x[100]);
  assign t[298] = (x[98]);
  assign t[299] = (x[87]);
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[106] & ~x[107] & ~x[108] & ~x[109]) | (~x[106] & x[107] & ~x[108] & ~x[109]) | (~x[106] & ~x[107] & x[108] & ~x[109]) | (~x[106] & ~x[107] & ~x[108] & x[109]) | (x[106] & x[107] & x[108] & ~x[109]) | (x[106] & x[107] & ~x[108] & x[109]) | (x[106] & ~x[107] & x[108] & x[109]) | (~x[106] & x[107] & x[108] & x[109]);
  assign t[301] = (x[108]);
  assign t[302] = (x[106]);
  assign t[303] = (x[101]);
  assign t[304] = (x[109]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[32] = t[48] ? x[31] : x[30];
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[44];
  assign t[38] = ~(t[107] & t[57]);
  assign t[39] = ~(t[108] & t[58]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[59] ? x[40] : x[39];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = ~(t[113] & t[74]);
  assign t[53] = t[103] ? x[57] : x[56];
  assign t[54] = ~(t[114] & t[75]);
  assign t[55] = ~(t[115] & t[76]);
  assign t[56] = t[103] ? x[66] : x[65];
  assign t[57] = ~(t[116]);
  assign t[58] = ~(t[116] & t[77]);
  assign t[59] = ~(t[25]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[117] & t[78]);
  assign t[61] = ~(t[118] & t[79]);
  assign t[62] = ~(t[119] & t[80]);
  assign t[63] = ~(t[120] & t[81]);
  assign t[64] = t[48] ? x[83] : x[82];
  assign t[65] = ~(t[82] & t[83]);
  assign t[66] = ~(t[121] & t[84]);
  assign t[67] = ~(t[122] & t[85]);
  assign t[68] = t[18] ? x[92] : x[91];
  assign t[69] = ~(t[86] & t[87]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[124]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[107]);
  assign t[78] = ~(t[126]);
  assign t[79] = ~(t[126] & t[91]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[114]);
  assign t[91] = ~(t[117]);
  assign t[92] = ~(t[119]);
  assign t[93] = ~(t[133]);
  assign t[94] = ~(t[133] & t[98]);
  assign t[95] = ~(t[121]);
  assign t[96] = ~(t[134]);
  assign t[97] = ~(t[134] & t[99]);
  assign t[98] = ~(t[128]);
  assign t[99] = ~(t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [124:0] x;
 output y;

 wire [466:0] t;
  assign t[0] = t[1] ? t[2] : t[212];
  assign t[100] = ~(t[147] & t[148]);
  assign t[101] = ~(t[234]);
  assign t[102] = ~(t[235]);
  assign t[103] = ~(t[149] | t[150]);
  assign t[104] = t[215] ? x[89] : x[88];
  assign t[105] = t[151] | t[152];
  assign t[106] = ~(t[236]);
  assign t[107] = ~(t[224] | t[225]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[238]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[153] | t[154]);
  assign t[111] = ~(t[140] | t[155]);
  assign t[112] = ~(t[156] | t[85]);
  assign t[113] = ~(t[239]);
  assign t[114] = ~(t[240]);
  assign t[115] = ~(t[157] | t[158]);
  assign t[116] = ~(t[159] | t[160]);
  assign t[117] = ~(t[241] | t[161]);
  assign t[118] = t[30] ? x[102] : x[101];
  assign t[119] = ~(t[162] & t[163]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[242]);
  assign t[121] = ~(t[243]);
  assign t[122] = ~(t[164] | t[165]);
  assign t[123] = ~(t[166] | t[167]);
  assign t[124] = ~(t[244] | t[168]);
  assign t[125] = t[30] ? x[112] : x[111];
  assign t[126] = ~(t[169] & t[170]);
  assign t[127] = ~(t[215]);
  assign t[128] = ~(t[171] & t[172]);
  assign t[129] = ~(t[173] & t[216]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[216] & t[174]);
  assign t[131] = ~(x[7] & t[175]);
  assign t[132] = ~(t[176] | t[142]);
  assign t[133] = ~(t[177] & t[178]);
  assign t[134] = t[213] ? t[130] : t[131];
  assign t[135] = ~(t[179]);
  assign t[136] = ~(t[82] | t[180]);
  assign t[137] = t[213] ? t[131] : t[181];
  assign t[138] = ~(t[245]);
  assign t[139] = ~(t[230] | t[231]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[82] | t[182]);
  assign t[141] = ~(t[31] & t[183]);
  assign t[142] = ~(t[127] | t[184]);
  assign t[143] = t[155] | t[135];
  assign t[144] = ~(t[246]);
  assign t[145] = ~(t[232] | t[233]);
  assign t[146] = ~(t[49]);
  assign t[147] = ~(t[151] | t[185]);
  assign t[148] = ~(t[140]);
  assign t[149] = ~(t[247]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[234] | t[235]);
  assign t[151] = ~(t[179] & t[133]);
  assign t[152] = ~(t[111] & t[186]);
  assign t[153] = ~(t[248]);
  assign t[154] = ~(t[237] | t[238]);
  assign t[155] = ~(t[82] | t[187]);
  assign t[156] = ~(t[127] | t[188]);
  assign t[157] = ~(t[249]);
  assign t[158] = ~(t[239] | t[240]);
  assign t[159] = ~(t[250]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[251]);
  assign t[161] = ~(t[189] | t[190]);
  assign t[162] = ~(t[156] | t[191]);
  assign t[163] = ~(t[155] | t[192]);
  assign t[164] = ~(t[252]);
  assign t[165] = ~(t[242] | t[243]);
  assign t[166] = ~(t[253]);
  assign t[167] = ~(t[254]);
  assign t[168] = ~(t[193] | t[194]);
  assign t[169] = ~(t[195] | t[196]);
  assign t[16] = ~(t[213] & t[214]);
  assign t[170] = ~(t[50] | t[197]);
  assign t[171] = ~(x[7] | t[214]);
  assign t[172] = ~(t[216]);
  assign t[173] = x[7] & t[214];
  assign t[174] = ~(x[7] | t[198]);
  assign t[175] = ~(t[214] | t[216]);
  assign t[176] = ~(t[127] | t[199]);
  assign t[177] = ~(t[214] | t[172]);
  assign t[178] = t[82] & t[213];
  assign t[179] = ~(t[200] & t[201]);
  assign t[17] = ~(t[215] & t[216]);
  assign t[180] = t[213] ? t[202] : t[181];
  assign t[181] = ~(t[174] & t[172]);
  assign t[182] = t[213] ? t[128] : t[129];
  assign t[183] = ~(t[203] & t[204]);
  assign t[184] = t[213] ? t[181] : t[131];
  assign t[185] = ~(t[205] & t[88]);
  assign t[186] = ~(t[51] | t[197]);
  assign t[187] = t[213] ? t[207] : t[206];
  assign t[188] = t[213] ? t[128] : t[206];
  assign t[189] = ~(t[255]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[250] | t[251]);
  assign t[191] = ~(t[82] | t[208]);
  assign t[192] = ~(t[170] & t[88]);
  assign t[193] = ~(t[256]);
  assign t[194] = ~(t[253] | t[254]);
  assign t[195] = ~(t[162] & t[209]);
  assign t[196] = ~(t[183] & t[88]);
  assign t[197] = ~(t[82] | t[210]);
  assign t[198] = ~(t[214]);
  assign t[199] = t[213] ? t[206] : t[128];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[127] | t[213]);
  assign t[201] = ~(t[130] & t[202]);
  assign t[202] = ~(x[7] & t[177]);
  assign t[203] = t[216] & t[200];
  assign t[204] = t[171] | t[173];
  assign t[205] = ~(t[142]);
  assign t[206] = ~(t[173] & t[172]);
  assign t[207] = ~(t[171] & t[216]);
  assign t[208] = t[213] ? t[181] : t[202];
  assign t[209] = ~(t[127] & t[211]);
  assign t[20] = t[30] ? x[9] : x[10];
  assign t[210] = t[213] ? t[206] : t[207];
  assign t[211] = ~(t[131] & t[130]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = (t[296]);
  assign t[252] = (t[297]);
  assign t[253] = (t[298]);
  assign t[254] = (t[299]);
  assign t[255] = (t[300]);
  assign t[256] = (t[301]);
  assign t[257] = t[302] ^ x[5];
  assign t[258] = t[303] ^ x[13];
  assign t[259] = t[304] ^ x[16];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[19];
  assign t[261] = t[306] ^ x[22];
  assign t[262] = t[307] ^ x[28];
  assign t[263] = t[308] ^ x[34];
  assign t[264] = t[309] ^ x[35];
  assign t[265] = t[310] ^ x[36];
  assign t[266] = t[311] ^ x[42];
  assign t[267] = t[312] ^ x[50];
  assign t[268] = t[313] ^ x[56];
  assign t[269] = t[314] ^ x[57];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[58];
  assign t[271] = t[316] ^ x[64];
  assign t[272] = t[317] ^ x[72];
  assign t[273] = t[318] ^ x[78];
  assign t[274] = t[319] ^ x[79];
  assign t[275] = t[320] ^ x[80];
  assign t[276] = t[321] ^ x[81];
  assign t[277] = t[322] ^ x[82];
  assign t[278] = t[323] ^ x[83];
  assign t[279] = t[324] ^ x[86];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[87];
  assign t[281] = t[326] ^ x[90];
  assign t[282] = t[327] ^ x[91];
  assign t[283] = t[328] ^ x[92];
  assign t[284] = t[329] ^ x[93];
  assign t[285] = t[330] ^ x[94];
  assign t[286] = t[331] ^ x[100];
  assign t[287] = t[332] ^ x[103];
  assign t[288] = t[333] ^ x[104];
  assign t[289] = t[334] ^ x[110];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[113];
  assign t[291] = t[336] ^ x[114];
  assign t[292] = t[337] ^ x[115];
  assign t[293] = t[338] ^ x[116];
  assign t[294] = t[339] ^ x[117];
  assign t[295] = t[340] ^ x[118];
  assign t[296] = t[341] ^ x[119];
  assign t[297] = t[342] ^ x[120];
  assign t[298] = t[343] ^ x[121];
  assign t[299] = t[344] ^ x[122];
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[345] ^ x[123];
  assign t[301] = t[346] ^ x[124];
  assign t[302] = (~t[347] & t[348]);
  assign t[303] = (~t[349] & t[350]);
  assign t[304] = (~t[351] & t[352]);
  assign t[305] = (~t[353] & t[354]);
  assign t[306] = (~t[355] & t[356]);
  assign t[307] = (~t[357] & t[358]);
  assign t[308] = (~t[359] & t[360]);
  assign t[309] = (~t[357] & t[361]);
  assign t[30] = ~(t[49]);
  assign t[310] = (~t[357] & t[362]);
  assign t[311] = (~t[363] & t[364]);
  assign t[312] = (~t[365] & t[366]);
  assign t[313] = (~t[367] & t[368]);
  assign t[314] = (~t[359] & t[369]);
  assign t[315] = (~t[359] & t[370]);
  assign t[316] = (~t[371] & t[372]);
  assign t[317] = (~t[373] & t[374]);
  assign t[318] = (~t[375] & t[376]);
  assign t[319] = (~t[357] & t[377]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (~t[363] & t[378]);
  assign t[321] = (~t[363] & t[379]);
  assign t[322] = (~t[365] & t[380]);
  assign t[323] = (~t[365] & t[381]);
  assign t[324] = (~t[367] & t[382]);
  assign t[325] = (~t[367] & t[383]);
  assign t[326] = (~t[359] & t[384]);
  assign t[327] = (~t[371] & t[385]);
  assign t[328] = (~t[371] & t[386]);
  assign t[329] = (~t[373] & t[387]);
  assign t[32] = ~(t[52] | t[53]);
  assign t[330] = (~t[373] & t[388]);
  assign t[331] = (~t[389] & t[390]);
  assign t[332] = (~t[375] & t[391]);
  assign t[333] = (~t[375] & t[392]);
  assign t[334] = (~t[393] & t[394]);
  assign t[335] = (~t[363] & t[395]);
  assign t[336] = (~t[365] & t[396]);
  assign t[337] = (~t[367] & t[397]);
  assign t[338] = (~t[371] & t[398]);
  assign t[339] = (~t[373] & t[399]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = (~t[389] & t[400]);
  assign t[341] = (~t[389] & t[401]);
  assign t[342] = (~t[375] & t[402]);
  assign t[343] = (~t[393] & t[403]);
  assign t[344] = (~t[393] & t[404]);
  assign t[345] = (~t[389] & t[405]);
  assign t[346] = (~t[393] & t[406]);
  assign t[347] = t[407] ^ x[4];
  assign t[348] = t[408] ^ x[5];
  assign t[349] = t[409] ^ x[12];
  assign t[34] = ~(t[217] | t[56]);
  assign t[350] = t[410] ^ x[13];
  assign t[351] = t[411] ^ x[15];
  assign t[352] = t[412] ^ x[16];
  assign t[353] = t[413] ^ x[18];
  assign t[354] = t[414] ^ x[19];
  assign t[355] = t[415] ^ x[21];
  assign t[356] = t[416] ^ x[22];
  assign t[357] = t[417] ^ x[27];
  assign t[358] = t[418] ^ x[28];
  assign t[359] = t[419] ^ x[33];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[420] ^ x[34];
  assign t[361] = t[421] ^ x[35];
  assign t[362] = t[422] ^ x[36];
  assign t[363] = t[423] ^ x[41];
  assign t[364] = t[424] ^ x[42];
  assign t[365] = t[425] ^ x[49];
  assign t[366] = t[426] ^ x[50];
  assign t[367] = t[427] ^ x[55];
  assign t[368] = t[428] ^ x[56];
  assign t[369] = t[429] ^ x[57];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[430] ^ x[58];
  assign t[371] = t[431] ^ x[63];
  assign t[372] = t[432] ^ x[64];
  assign t[373] = t[433] ^ x[71];
  assign t[374] = t[434] ^ x[72];
  assign t[375] = t[435] ^ x[77];
  assign t[376] = t[436] ^ x[78];
  assign t[377] = t[437] ^ x[79];
  assign t[378] = t[438] ^ x[80];
  assign t[379] = t[439] ^ x[81];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[440] ^ x[82];
  assign t[381] = t[441] ^ x[83];
  assign t[382] = t[442] ^ x[86];
  assign t[383] = t[443] ^ x[87];
  assign t[384] = t[444] ^ x[90];
  assign t[385] = t[445] ^ x[91];
  assign t[386] = t[446] ^ x[92];
  assign t[387] = t[447] ^ x[93];
  assign t[388] = t[448] ^ x[94];
  assign t[389] = t[449] ^ x[99];
  assign t[38] = ~(t[45] ^ t[63]);
  assign t[390] = t[450] ^ x[100];
  assign t[391] = t[451] ^ x[103];
  assign t[392] = t[452] ^ x[104];
  assign t[393] = t[453] ^ x[109];
  assign t[394] = t[454] ^ x[110];
  assign t[395] = t[455] ^ x[113];
  assign t[396] = t[456] ^ x[114];
  assign t[397] = t[457] ^ x[115];
  assign t[398] = t[458] ^ x[116];
  assign t[399] = t[459] ^ x[117];
  assign t[39] = ~(t[64] | t[65]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[460] ^ x[118];
  assign t[401] = t[461] ^ x[119];
  assign t[402] = t[462] ^ x[120];
  assign t[403] = t[463] ^ x[121];
  assign t[404] = t[464] ^ x[122];
  assign t[405] = t[465] ^ x[123];
  assign t[406] = t[466] ^ x[124];
  assign t[407] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[408] = (x[0]);
  assign t[409] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[40] = ~(t[39] ^ t[66]);
  assign t[410] = (x[11]);
  assign t[411] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[412] = (x[14]);
  assign t[413] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[414] = (x[17]);
  assign t[415] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[416] = (x[20]);
  assign t[417] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[418] = (x[24]);
  assign t[419] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[420] = (x[30]);
  assign t[421] = (x[25]);
  assign t[422] = (x[26]);
  assign t[423] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[424] = (x[38]);
  assign t[425] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[426] = (x[46]);
  assign t[427] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[428] = (x[52]);
  assign t[429] = (x[31]);
  assign t[42] = ~(t[218] | t[69]);
  assign t[430] = (x[32]);
  assign t[431] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[432] = (x[60]);
  assign t[433] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[434] = (x[68]);
  assign t[435] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[436] = (x[74]);
  assign t[437] = (x[23]);
  assign t[438] = (x[39]);
  assign t[439] = (x[40]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (x[47]);
  assign t[441] = (x[48]);
  assign t[442] = (x[53]);
  assign t[443] = (x[54]);
  assign t[444] = (x[29]);
  assign t[445] = (x[61]);
  assign t[446] = (x[62]);
  assign t[447] = (x[69]);
  assign t[448] = (x[70]);
  assign t[449] = (x[95] & ~x[96] & ~x[97] & ~x[98]) | (~x[95] & x[96] & ~x[97] & ~x[98]) | (~x[95] & ~x[96] & x[97] & ~x[98]) | (~x[95] & ~x[96] & ~x[97] & x[98]) | (x[95] & x[96] & x[97] & ~x[98]) | (x[95] & x[96] & ~x[97] & x[98]) | (x[95] & ~x[96] & x[97] & x[98]) | (~x[95] & x[96] & x[97] & x[98]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (x[96]);
  assign t[451] = (x[75]);
  assign t[452] = (x[76]);
  assign t[453] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[454] = (x[106]);
  assign t[455] = (x[37]);
  assign t[456] = (x[45]);
  assign t[457] = (x[51]);
  assign t[458] = (x[59]);
  assign t[459] = (x[67]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = (x[97]);
  assign t[461] = (x[98]);
  assign t[462] = (x[73]);
  assign t[463] = (x[107]);
  assign t[464] = (x[108]);
  assign t[465] = (x[95]);
  assign t[466] = (x[105]);
  assign t[46] = ~(t[76] ^ t[77]);
  assign t[47] = ~(t[78] | t[79]);
  assign t[48] = ~(t[80] ^ t[81]);
  assign t[49] = ~(t[215]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[82] | t[83]);
  assign t[51] = ~(t[82] | t[84]);
  assign t[52] = t[85] | t[86];
  assign t[53] = ~(t[87] & t[88]);
  assign t[54] = ~(t[219]);
  assign t[55] = ~(t[220]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[221] | t[93]);
  assign t[59] = t[215] ? x[44] : x[43];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[222] | t[98]);
  assign t[63] = ~(t[99] ^ t[100]);
  assign t[64] = ~(t[101] | t[102]);
  assign t[65] = ~(t[223] | t[103]);
  assign t[66] = ~(t[104] ^ t[105]);
  assign t[67] = ~(t[224]);
  assign t[68] = ~(t[225]);
  assign t[69] = ~(t[106] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[226] | t[110]);
  assign t[72] = t[30] ? x[66] : x[65];
  assign t[73] = ~(t[111] & t[112]);
  assign t[74] = ~(t[113] | t[114]);
  assign t[75] = ~(t[227] | t[115]);
  assign t[76] = ~(t[116] | t[117]);
  assign t[77] = ~(t[118] ^ t[119]);
  assign t[78] = ~(t[120] | t[121]);
  assign t[79] = ~(t[228] | t[122]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[123] | t[124]);
  assign t[81] = ~(t[125] ^ t[126]);
  assign t[82] = ~(t[127]);
  assign t[83] = t[213] ? t[129] : t[128];
  assign t[84] = t[213] ? t[131] : t[130];
  assign t[85] = ~(t[132] & t[133]);
  assign t[86] = ~(t[82] | t[134]);
  assign t[87] = ~(t[135] | t[136]);
  assign t[88] = t[127] | t[137];
  assign t[89] = ~(t[229]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[219] | t[220]);
  assign t[91] = ~(t[230]);
  assign t[92] = ~(t[231]);
  assign t[93] = ~(t[138] | t[139]);
  assign t[94] = ~(t[140] | t[141]);
  assign t[95] = ~(t[142] | t[143]);
  assign t[96] = ~(t[232]);
  assign t[97] = ~(t[233]);
  assign t[98] = ~(t[144] | t[145]);
  assign t[99] = t[146] ? x[85] : x[84];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [163:0] x;
 output y;

 wire [629:0] t;
  assign t[0] = t[1] ? t[2] : t[382];
  assign t[100] = ~(t[404]);
  assign t[101] = ~(t[393] | t[394]);
  assign t[102] = ~(t[405]);
  assign t[103] = ~(t[406]);
  assign t[104] = ~(t[138] | t[139]);
  assign t[105] = ~(t[86] | t[140]);
  assign t[106] = ~(t[141] & t[142]);
  assign t[107] = ~(t[407]);
  assign t[108] = ~(t[408]);
  assign t[109] = ~(t[143] | t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[145] ? x[94] : x[93];
  assign t[111] = t[146] | t[147];
  assign t[112] = ~(t[409]);
  assign t[113] = ~(t[410]);
  assign t[114] = ~(t[148] | t[149]);
  assign t[115] = ~(t[150] | t[151]);
  assign t[116] = ~(t[411] | t[152]);
  assign t[117] = t[145] ? x[104] : x[103];
  assign t[118] = ~(t[153] & t[154]);
  assign t[119] = ~(t[385]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[155] & t[83]);
  assign t[121] = ~(t[156] & t[386]);
  assign t[122] = ~(t[119] | t[157]);
  assign t[123] = ~(t[79] | t[158]);
  assign t[124] = ~(t[159] & t[160]);
  assign t[125] = ~(t[161] & t[162]);
  assign t[126] = ~(t[163] | t[164]);
  assign t[127] = ~(t[165] | t[166]);
  assign t[128] = ~(t[412]);
  assign t[129] = ~(t[399] | t[400]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[163] | t[167]);
  assign t[131] = ~(t[168] | t[169]);
  assign t[132] = ~(t[413]);
  assign t[133] = ~(t[401] | t[402]);
  assign t[134] = ~(t[414]);
  assign t[135] = ~(t[415]);
  assign t[136] = ~(t[170] | t[171]);
  assign t[137] = ~(t[172] | t[166]);
  assign t[138] = ~(t[416]);
  assign t[139] = ~(t[405] | t[406]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[147] | t[164];
  assign t[141] = t[386] & t[161];
  assign t[142] = t[155] | t[156];
  assign t[143] = ~(t[417]);
  assign t[144] = ~(t[407] | t[408]);
  assign t[145] = ~(t[48]);
  assign t[146] = ~(t[173] & t[32]);
  assign t[147] = ~(t[79] | t[174]);
  assign t[148] = ~(t[418]);
  assign t[149] = ~(t[409] | t[410]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[419]);
  assign t[151] = ~(t[420]);
  assign t[152] = ~(t[175] | t[176]);
  assign t[153] = ~(t[49]);
  assign t[154] = ~(t[177] | t[147]);
  assign t[155] = ~(x[7] | t[384]);
  assign t[156] = x[7] & t[384];
  assign t[157] = t[383] ? t[120] : t[178];
  assign t[158] = t[383] ? t[180] : t[179];
  assign t[159] = ~(x[7] & t[181]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[386] & t[182]);
  assign t[161] = ~(t[119] | t[383]);
  assign t[162] = ~(t[160] & t[179]);
  assign t[163] = ~(t[79] | t[183]);
  assign t[164] = ~(t[79] | t[184]);
  assign t[165] = ~(t[79] | t[185]);
  assign t[166] = ~(t[79] | t[186]);
  assign t[167] = ~(t[187] & t[106]);
  assign t[168] = ~(t[119] | t[188]);
  assign t[169] = t[164] | t[189];
  assign t[16] = ~(t[383] & t[384]);
  assign t[170] = ~(t[421]);
  assign t[171] = ~(t[414] | t[415]);
  assign t[172] = ~(t[79] | t[190]);
  assign t[173] = ~(t[191] | t[168]);
  assign t[174] = t[383] ? t[160] : t[159];
  assign t[175] = ~(t[422]);
  assign t[176] = ~(t[419] | t[420]);
  assign t[177] = ~(t[137]);
  assign t[178] = ~(t[156] & t[83]);
  assign t[179] = ~(x[7] & t[51]);
  assign t[17] = ~(t[385] & t[386]);
  assign t[180] = ~(t[182] & t[83]);
  assign t[181] = ~(t[384] | t[386]);
  assign t[182] = ~(x[7] | t[192]);
  assign t[183] = t[383] ? t[120] : t[121];
  assign t[184] = t[383] ? t[193] : t[178];
  assign t[185] = t[383] ? t[159] : t[160];
  assign t[186] = t[383] ? t[178] : t[193];
  assign t[187] = ~(t[49] | t[165]);
  assign t[188] = t[383] ? t[180] : t[159];
  assign t[189] = ~(t[125]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = t[383] ? t[179] : t[180];
  assign t[191] = ~(t[119] | t[194]);
  assign t[192] = ~(t[384]);
  assign t[193] = ~(t[155] & t[386]);
  assign t[194] = t[383] ? t[178] : t[120];
  assign t[195] = t[1] ? t[196] : t[423];
  assign t[196] = x[6] ? t[198] : t[197];
  assign t[197] = x[7] ? t[200] : t[199];
  assign t[198] = t[201] ^ x[117];
  assign t[199] = t[202] ^ t[203];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[204] ^ t[205]);
  assign t[201] = x[118] ^ x[119];
  assign t[202] = t[30] ? x[118] : x[119];
  assign t[203] = ~(t[206] ^ t[207]);
  assign t[204] = x[7] ? t[209] : t[208];
  assign t[205] = ~(t[210] ^ t[211]);
  assign t[206] = x[7] ? t[213] : t[212];
  assign t[207] = ~(t[214] ^ t[215]);
  assign t[208] = ~(t[216] & t[217]);
  assign t[209] = t[218] ^ t[208];
  assign t[20] = t[30] ? x[9] : x[10];
  assign t[210] = x[7] ? t[220] : t[219];
  assign t[211] = x[7] ? t[222] : t[221];
  assign t[212] = ~(t[223] & t[224]);
  assign t[213] = t[225] ^ t[226];
  assign t[214] = x[7] ? t[228] : t[227];
  assign t[215] = x[7] ? t[230] : t[229];
  assign t[216] = ~(t[389] & t[54]);
  assign t[217] = ~(t[398] & t[231]);
  assign t[218] = t[385] ? x[121] : x[120];
  assign t[219] = ~(t[232] & t[233]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = t[234] ^ t[235];
  assign t[221] = ~(t[236] & t[237]);
  assign t[222] = t[238] ^ t[229];
  assign t[223] = ~(t[393] & t[66]);
  assign t[224] = ~(t[404] & t[239]);
  assign t[225] = t[30] ? x[123] : x[122];
  assign t[226] = ~(t[240] & t[241]);
  assign t[227] = ~(t[242] & t[243]);
  assign t[228] = t[244] ^ t[245];
  assign t[229] = ~(t[246] & t[247]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = t[248] ^ t[227];
  assign t[231] = ~(t[390] & t[53]);
  assign t[232] = ~(t[401] & t[94]);
  assign t[233] = ~(t[413] & t[249]);
  assign t[234] = t[385] ? x[125] : x[124];
  assign t[235] = ~(t[250] & t[251]);
  assign t[236] = ~(t[399] & t[89]);
  assign t[237] = ~(t[412] & t[252]);
  assign t[238] = t[253] ? x[127] : x[126];
  assign t[239] = ~(t[394] & t[65]);
  assign t[23] = ~(t[22] ^ t[35]);
  assign t[240] = ~(t[405] & t[103]);
  assign t[241] = ~(t[416] & t[254]);
  assign t[242] = ~(t[409] & t[113]);
  assign t[243] = ~(t[418] & t[255]);
  assign t[244] = t[145] ? x[129] : x[128];
  assign t[245] = ~(t[256] & t[257]);
  assign t[246] = ~(t[407] & t[108]);
  assign t[247] = ~(t[417] & t[258]);
  assign t[248] = t[145] ? x[131] : x[130];
  assign t[249] = ~(t[402] & t[93]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = ~(t[414] & t[135]);
  assign t[251] = ~(t[421] & t[259]);
  assign t[252] = ~(t[400] & t[88]);
  assign t[253] = ~(t[48]);
  assign t[254] = ~(t[406] & t[102]);
  assign t[255] = ~(t[410] & t[112]);
  assign t[256] = ~(t[419] & t[151]);
  assign t[257] = ~(t[422] & t[260]);
  assign t[258] = ~(t[408] & t[107]);
  assign t[259] = ~(t[415] & t[134]);
  assign t[25] = x[7] ? t[39] : t[38];
  assign t[260] = ~(t[420] & t[150]);
  assign t[261] = t[1] ? t[262] : t[424];
  assign t[262] = x[6] ? t[264] : t[263];
  assign t[263] = x[7] ? t[266] : t[265];
  assign t[264] = t[267] ^ x[133];
  assign t[265] = t[268] ^ t[269];
  assign t[266] = ~(t[270] ^ t[271]);
  assign t[267] = x[134] ^ x[135];
  assign t[268] = t[30] ? x[134] : x[135];
  assign t[269] = ~(t[272] ^ t[273]);
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = x[7] ? t[275] : t[274];
  assign t[271] = ~(t[276] ^ t[277]);
  assign t[272] = x[7] ? t[279] : t[278];
  assign t[273] = ~(t[280] ^ t[281]);
  assign t[274] = ~(t[282] & t[283]);
  assign t[275] = t[284] ^ t[274];
  assign t[276] = x[7] ? t[286] : t[285];
  assign t[277] = x[7] ? t[288] : t[287];
  assign t[278] = ~(t[289] & t[290]);
  assign t[279] = t[291] ^ t[292];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = x[7] ? t[294] : t[293];
  assign t[281] = x[7] ? t[296] : t[295];
  assign t[282] = ~(t[54] & t[84]);
  assign t[283] = ~(t[297] & t[387]);
  assign t[284] = t[385] ? x[137] : x[136];
  assign t[285] = ~(t[298] & t[299]);
  assign t[286] = t[300] ^ t[301];
  assign t[287] = ~(t[302] & t[303]);
  assign t[288] = t[304] ^ t[293];
  assign t[289] = ~(t[66] & t[100]);
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = ~(t[305] & t[388]);
  assign t[291] = t[30] ? x[139] : x[138];
  assign t[292] = ~(t[306] & t[307]);
  assign t[293] = ~(t[308] & t[309]);
  assign t[294] = t[310] ^ t[295];
  assign t[295] = ~(t[311] & t[312]);
  assign t[296] = t[313] ^ t[314];
  assign t[297] = ~(t[315] & t[53]);
  assign t[298] = ~(t[94] & t[132]);
  assign t[299] = ~(t[316] & t[392]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[385] ? x[141] : x[140];
  assign t[301] = ~(t[317] & t[318]);
  assign t[302] = ~(t[89] & t[128]);
  assign t[303] = ~(t[319] & t[391]);
  assign t[304] = t[30] ? x[143] : x[142];
  assign t[305] = ~(t[320] & t[65]);
  assign t[306] = ~(t[103] & t[138]);
  assign t[307] = ~(t[321] & t[395]);
  assign t[308] = ~(t[108] & t[143]);
  assign t[309] = ~(t[322] & t[396]);
  assign t[30] = ~(t[48]);
  assign t[310] = t[145] ? x[145] : x[144];
  assign t[311] = ~(t[113] & t[148]);
  assign t[312] = ~(t[323] & t[397]);
  assign t[313] = t[145] ? x[147] : x[146];
  assign t[314] = ~(t[324] & t[325]);
  assign t[315] = ~(t[398] & t[390]);
  assign t[316] = ~(t[326] & t[93]);
  assign t[317] = ~(t[135] & t[170]);
  assign t[318] = ~(t[327] & t[403]);
  assign t[319] = ~(t[328] & t[88]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = ~(t[404] & t[394]);
  assign t[321] = ~(t[329] & t[102]);
  assign t[322] = ~(t[330] & t[107]);
  assign t[323] = ~(t[331] & t[112]);
  assign t[324] = ~(t[151] & t[175]);
  assign t[325] = ~(t[332] & t[411]);
  assign t[326] = ~(t[413] & t[402]);
  assign t[327] = ~(t[333] & t[134]);
  assign t[328] = ~(t[412] & t[400]);
  assign t[329] = ~(t[416] & t[406]);
  assign t[32] = ~(t[51] & t[52]);
  assign t[330] = ~(t[417] & t[408]);
  assign t[331] = ~(t[418] & t[410]);
  assign t[332] = ~(t[334] & t[150]);
  assign t[333] = ~(t[421] & t[415]);
  assign t[334] = ~(t[422] & t[420]);
  assign t[335] = t[1] ? t[336] : t[425];
  assign t[336] = x[6] ? t[338] : t[337];
  assign t[337] = x[7] ? t[340] : t[339];
  assign t[338] = t[341] ^ x[149];
  assign t[339] = t[342] ^ t[343];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = ~(t[344] ^ t[345]);
  assign t[341] = x[150] ^ x[151];
  assign t[342] = t[30] ? x[150] : x[151];
  assign t[343] = ~(t[346] ^ t[347]);
  assign t[344] = x[7] ? t[349] : t[348];
  assign t[345] = ~(t[350] ^ t[351]);
  assign t[346] = x[7] ? t[353] : t[352];
  assign t[347] = ~(t[354] ^ t[355]);
  assign t[348] = ~(t[282] & t[356]);
  assign t[349] = t[357] ^ t[348];
  assign t[34] = ~(t[387] | t[55]);
  assign t[350] = x[7] ? t[359] : t[358];
  assign t[351] = x[7] ? t[361] : t[360];
  assign t[352] = ~(t[289] & t[362]);
  assign t[353] = t[363] ^ t[364];
  assign t[354] = x[7] ? t[366] : t[365];
  assign t[355] = x[7] ? t[368] : t[367];
  assign t[356] = t[33] | t[387];
  assign t[357] = t[385] ? x[153] : x[152];
  assign t[358] = ~(t[298] & t[369]);
  assign t[359] = t[370] ^ t[371];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = ~(t[302] & t[372]);
  assign t[361] = t[373] ^ t[365];
  assign t[362] = t[40] | t[388];
  assign t[363] = t[30] ? x[155] : x[154];
  assign t[364] = ~(t[306] & t[374]);
  assign t[365] = ~(t[308] & t[375]);
  assign t[366] = t[376] ^ t[367];
  assign t[367] = ~(t[311] & t[377]);
  assign t[368] = t[378] ^ t[379];
  assign t[369] = t[61] | t[392];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[385] ? x[157] : x[156];
  assign t[371] = ~(t[317] & t[380]);
  assign t[372] = t[58] | t[391];
  assign t[373] = t[145] ? x[159] : x[158];
  assign t[374] = t[68] | t[395];
  assign t[375] = t[72] | t[396];
  assign t[376] = t[145] ? x[161] : x[160];
  assign t[377] = t[75] | t[397];
  assign t[378] = t[145] ? x[163] : x[162];
  assign t[379] = ~(t[324] & t[381]);
  assign t[37] = ~(t[44] ^ t[60]);
  assign t[380] = t[96] | t[403];
  assign t[381] = t[115] | t[411];
  assign t[382] = (t[426]);
  assign t[383] = (t[427]);
  assign t[384] = (t[428]);
  assign t[385] = (t[429]);
  assign t[386] = (t[430]);
  assign t[387] = (t[431]);
  assign t[388] = (t[432]);
  assign t[389] = (t[433]);
  assign t[38] = ~(t[61] | t[62]);
  assign t[390] = (t[434]);
  assign t[391] = (t[435]);
  assign t[392] = (t[436]);
  assign t[393] = (t[437]);
  assign t[394] = (t[438]);
  assign t[395] = (t[439]);
  assign t[396] = (t[440]);
  assign t[397] = (t[441]);
  assign t[398] = (t[442]);
  assign t[399] = (t[443]);
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (t[444]);
  assign t[401] = (t[445]);
  assign t[402] = (t[446]);
  assign t[403] = (t[447]);
  assign t[404] = (t[448]);
  assign t[405] = (t[449]);
  assign t[406] = (t[450]);
  assign t[407] = (t[451]);
  assign t[408] = (t[452]);
  assign t[409] = (t[453]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (t[454]);
  assign t[411] = (t[455]);
  assign t[412] = (t[456]);
  assign t[413] = (t[457]);
  assign t[414] = (t[458]);
  assign t[415] = (t[459]);
  assign t[416] = (t[460]);
  assign t[417] = (t[461]);
  assign t[418] = (t[462]);
  assign t[419] = (t[463]);
  assign t[41] = ~(t[388] | t[67]);
  assign t[420] = (t[464]);
  assign t[421] = (t[465]);
  assign t[422] = (t[466]);
  assign t[423] = (t[467]);
  assign t[424] = (t[468]);
  assign t[425] = (t[469]);
  assign t[426] = t[470] ^ x[5];
  assign t[427] = t[471] ^ x[13];
  assign t[428] = t[472] ^ x[16];
  assign t[429] = t[473] ^ x[19];
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = t[474] ^ x[22];
  assign t[431] = t[475] ^ x[28];
  assign t[432] = t[476] ^ x[34];
  assign t[433] = t[477] ^ x[35];
  assign t[434] = t[478] ^ x[36];
  assign t[435] = t[479] ^ x[44];
  assign t[436] = t[480] ^ x[50];
  assign t[437] = t[481] ^ x[51];
  assign t[438] = t[482] ^ x[52];
  assign t[439] = t[483] ^ x[58];
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = t[484] ^ x[66];
  assign t[441] = t[485] ^ x[72];
  assign t[442] = t[486] ^ x[73];
  assign t[443] = t[487] ^ x[74];
  assign t[444] = t[488] ^ x[75];
  assign t[445] = t[489] ^ x[78];
  assign t[446] = t[490] ^ x[79];
  assign t[447] = t[491] ^ x[85];
  assign t[448] = t[492] ^ x[88];
  assign t[449] = t[493] ^ x[89];
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = t[494] ^ x[90];
  assign t[451] = t[495] ^ x[91];
  assign t[452] = t[496] ^ x[92];
  assign t[453] = t[497] ^ x[95];
  assign t[454] = t[498] ^ x[96];
  assign t[455] = t[499] ^ x[102];
  assign t[456] = t[500] ^ x[105];
  assign t[457] = t[501] ^ x[106];
  assign t[458] = t[502] ^ x[107];
  assign t[459] = t[503] ^ x[108];
  assign t[45] = ~(t[46] ^ t[74]);
  assign t[460] = t[504] ^ x[109];
  assign t[461] = t[505] ^ x[110];
  assign t[462] = t[506] ^ x[111];
  assign t[463] = t[507] ^ x[112];
  assign t[464] = t[508] ^ x[113];
  assign t[465] = t[509] ^ x[114];
  assign t[466] = t[510] ^ x[115];
  assign t[467] = t[511] ^ x[116];
  assign t[468] = t[512] ^ x[132];
  assign t[469] = t[513] ^ x[148];
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = (~t[514] & t[515]);
  assign t[471] = (~t[516] & t[517]);
  assign t[472] = (~t[518] & t[519]);
  assign t[473] = (~t[520] & t[521]);
  assign t[474] = (~t[522] & t[523]);
  assign t[475] = (~t[524] & t[525]);
  assign t[476] = (~t[526] & t[527]);
  assign t[477] = (~t[524] & t[528]);
  assign t[478] = (~t[524] & t[529]);
  assign t[479] = (~t[530] & t[531]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (~t[532] & t[533]);
  assign t[481] = (~t[526] & t[534]);
  assign t[482] = (~t[526] & t[535]);
  assign t[483] = (~t[536] & t[537]);
  assign t[484] = (~t[538] & t[539]);
  assign t[485] = (~t[540] & t[541]);
  assign t[486] = (~t[524] & t[542]);
  assign t[487] = (~t[530] & t[543]);
  assign t[488] = (~t[530] & t[544]);
  assign t[489] = (~t[532] & t[545]);
  assign t[48] = ~(t[385]);
  assign t[490] = (~t[532] & t[546]);
  assign t[491] = (~t[547] & t[548]);
  assign t[492] = (~t[526] & t[549]);
  assign t[493] = (~t[536] & t[550]);
  assign t[494] = (~t[536] & t[551]);
  assign t[495] = (~t[538] & t[552]);
  assign t[496] = (~t[538] & t[553]);
  assign t[497] = (~t[540] & t[554]);
  assign t[498] = (~t[540] & t[555]);
  assign t[499] = (~t[556] & t[557]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[530] & t[558]);
  assign t[501] = (~t[532] & t[559]);
  assign t[502] = (~t[547] & t[560]);
  assign t[503] = (~t[547] & t[561]);
  assign t[504] = (~t[536] & t[562]);
  assign t[505] = (~t[538] & t[563]);
  assign t[506] = (~t[540] & t[564]);
  assign t[507] = (~t[556] & t[565]);
  assign t[508] = (~t[556] & t[566]);
  assign t[509] = (~t[547] & t[567]);
  assign t[50] = ~(t[81] & t[82]);
  assign t[510] = (~t[556] & t[568]);
  assign t[511] = (~t[514] & t[569]);
  assign t[512] = (~t[514] & t[570]);
  assign t[513] = (~t[514] & t[571]);
  assign t[514] = t[572] ^ x[4];
  assign t[515] = t[573] ^ x[5];
  assign t[516] = t[574] ^ x[12];
  assign t[517] = t[575] ^ x[13];
  assign t[518] = t[576] ^ x[15];
  assign t[519] = t[577] ^ x[16];
  assign t[51] = ~(t[384] | t[83]);
  assign t[520] = t[578] ^ x[18];
  assign t[521] = t[579] ^ x[19];
  assign t[522] = t[580] ^ x[21];
  assign t[523] = t[581] ^ x[22];
  assign t[524] = t[582] ^ x[27];
  assign t[525] = t[583] ^ x[28];
  assign t[526] = t[584] ^ x[33];
  assign t[527] = t[585] ^ x[34];
  assign t[528] = t[586] ^ x[35];
  assign t[529] = t[587] ^ x[36];
  assign t[52] = t[79] & t[383];
  assign t[530] = t[588] ^ x[43];
  assign t[531] = t[589] ^ x[44];
  assign t[532] = t[590] ^ x[49];
  assign t[533] = t[591] ^ x[50];
  assign t[534] = t[592] ^ x[51];
  assign t[535] = t[593] ^ x[52];
  assign t[536] = t[594] ^ x[57];
  assign t[537] = t[595] ^ x[58];
  assign t[538] = t[596] ^ x[65];
  assign t[539] = t[597] ^ x[66];
  assign t[53] = ~(t[389]);
  assign t[540] = t[598] ^ x[71];
  assign t[541] = t[599] ^ x[72];
  assign t[542] = t[600] ^ x[73];
  assign t[543] = t[601] ^ x[74];
  assign t[544] = t[602] ^ x[75];
  assign t[545] = t[603] ^ x[78];
  assign t[546] = t[604] ^ x[79];
  assign t[547] = t[605] ^ x[84];
  assign t[548] = t[606] ^ x[85];
  assign t[549] = t[607] ^ x[88];
  assign t[54] = ~(t[390]);
  assign t[550] = t[608] ^ x[89];
  assign t[551] = t[609] ^ x[90];
  assign t[552] = t[610] ^ x[91];
  assign t[553] = t[611] ^ x[92];
  assign t[554] = t[612] ^ x[95];
  assign t[555] = t[613] ^ x[96];
  assign t[556] = t[614] ^ x[101];
  assign t[557] = t[615] ^ x[102];
  assign t[558] = t[616] ^ x[105];
  assign t[559] = t[617] ^ x[106];
  assign t[55] = ~(t[84] | t[85]);
  assign t[560] = t[618] ^ x[107];
  assign t[561] = t[619] ^ x[108];
  assign t[562] = t[620] ^ x[109];
  assign t[563] = t[621] ^ x[110];
  assign t[564] = t[622] ^ x[111];
  assign t[565] = t[623] ^ x[112];
  assign t[566] = t[624] ^ x[113];
  assign t[567] = t[625] ^ x[114];
  assign t[568] = t[626] ^ x[115];
  assign t[569] = t[627] ^ x[116];
  assign t[56] = t[385] ? x[38] : x[37];
  assign t[570] = t[628] ^ x[132];
  assign t[571] = t[629] ^ x[148];
  assign t[572] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[573] = (x[0]);
  assign t[574] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[575] = (x[11]);
  assign t[576] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[577] = (x[14]);
  assign t[578] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[579] = (x[17]);
  assign t[57] = t[86] | t[87];
  assign t[580] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[581] = (x[20]);
  assign t[582] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[583] = (x[24]);
  assign t[584] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[585] = (x[30]);
  assign t[586] = (x[25]);
  assign t[587] = (x[26]);
  assign t[588] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[589] = (x[40]);
  assign t[58] = ~(t[88] | t[89]);
  assign t[590] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[591] = (x[46]);
  assign t[592] = (x[31]);
  assign t[593] = (x[32]);
  assign t[594] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[595] = (x[54]);
  assign t[596] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[597] = (x[62]);
  assign t[598] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[599] = (x[68]);
  assign t[59] = ~(t[391] | t[90]);
  assign t[5] = t[9] ^ x[8];
  assign t[600] = (x[23]);
  assign t[601] = (x[41]);
  assign t[602] = (x[42]);
  assign t[603] = (x[47]);
  assign t[604] = (x[48]);
  assign t[605] = (x[80] & ~x[81] & ~x[82] & ~x[83]) | (~x[80] & x[81] & ~x[82] & ~x[83]) | (~x[80] & ~x[81] & x[82] & ~x[83]) | (~x[80] & ~x[81] & ~x[82] & x[83]) | (x[80] & x[81] & x[82] & ~x[83]) | (x[80] & x[81] & ~x[82] & x[83]) | (x[80] & ~x[81] & x[82] & x[83]) | (~x[80] & x[81] & x[82] & x[83]);
  assign t[606] = (x[81]);
  assign t[607] = (x[29]);
  assign t[608] = (x[55]);
  assign t[609] = (x[56]);
  assign t[60] = ~(t[91] ^ t[92]);
  assign t[610] = (x[63]);
  assign t[611] = (x[64]);
  assign t[612] = (x[69]);
  assign t[613] = (x[70]);
  assign t[614] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[615] = (x[98]);
  assign t[616] = (x[39]);
  assign t[617] = (x[45]);
  assign t[618] = (x[82]);
  assign t[619] = (x[83]);
  assign t[61] = ~(t[93] | t[94]);
  assign t[620] = (x[53]);
  assign t[621] = (x[61]);
  assign t[622] = (x[67]);
  assign t[623] = (x[99]);
  assign t[624] = (x[100]);
  assign t[625] = (x[80]);
  assign t[626] = (x[97]);
  assign t[627] = (x[1]);
  assign t[628] = (x[2]);
  assign t[629] = (x[3]);
  assign t[62] = ~(t[392] | t[95]);
  assign t[63] = ~(t[96] | t[97]);
  assign t[64] = ~(t[98] ^ t[99]);
  assign t[65] = ~(t[393]);
  assign t[66] = ~(t[394]);
  assign t[67] = ~(t[100] | t[101]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[395] | t[104]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[30] ? x[60] : x[59];
  assign t[71] = ~(t[105] & t[106]);
  assign t[72] = ~(t[107] | t[108]);
  assign t[73] = ~(t[396] | t[109]);
  assign t[74] = ~(t[110] ^ t[111]);
  assign t[75] = ~(t[112] | t[113]);
  assign t[76] = ~(t[397] | t[114]);
  assign t[77] = ~(t[115] | t[116]);
  assign t[78] = ~(t[117] ^ t[118]);
  assign t[79] = ~(t[119]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[383] ? t[121] : t[120];
  assign t[81] = ~(t[122] | t[123]);
  assign t[82] = ~(t[119] & t[124]);
  assign t[83] = ~(t[386]);
  assign t[84] = ~(t[398]);
  assign t[85] = ~(t[389] | t[390]);
  assign t[86] = ~(t[125] & t[32]);
  assign t[87] = ~(t[126] & t[127]);
  assign t[88] = ~(t[399]);
  assign t[89] = ~(t[400]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[128] | t[129]);
  assign t[91] = t[385] ? x[77] : x[76];
  assign t[92] = ~(t[130] & t[131]);
  assign t[93] = ~(t[401]);
  assign t[94] = ~(t[402]);
  assign t[95] = ~(t[132] | t[133]);
  assign t[96] = ~(t[134] | t[135]);
  assign t[97] = ~(t[403] | t[136]);
  assign t[98] = t[385] ? x[87] : x[86];
  assign t[99] = ~(t[130] & t[137]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[195] & ~t[261] & ~t[335]) | (~t[0] & t[195] & ~t[261] & ~t[335]) | (~t[0] & ~t[195] & t[261] & ~t[335]) | (~t[0] & ~t[195] & ~t[261] & t[335]) | (t[0] & t[195] & t[261] & ~t[335]) | (t[0] & t[195] & ~t[261] & t[335]) | (t[0] & ~t[195] & t[261] & t[335]) | (~t[0] & t[195] & t[261] & t[335]);
endmodule

module R2ind151(x, y);
 input [115:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = t[1] ? t[2] : t[102];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = t[184] ^ x[5];
  assign t[144] = t[185] ^ x[13];
  assign t[145] = t[186] ^ x[16];
  assign t[146] = t[187] ^ x[19];
  assign t[147] = t[188] ^ x[22];
  assign t[148] = t[189] ^ x[28];
  assign t[149] = t[190] ^ x[36];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[39];
  assign t[151] = t[192] ^ x[40];
  assign t[152] = t[193] ^ x[46];
  assign t[153] = t[194] ^ x[54];
  assign t[154] = t[195] ^ x[57];
  assign t[155] = t[196] ^ x[58];
  assign t[156] = t[197] ^ x[64];
  assign t[157] = t[198] ^ x[70];
  assign t[158] = t[199] ^ x[78];
  assign t[159] = t[200] ^ x[81];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[82];
  assign t[161] = t[202] ^ x[83];
  assign t[162] = t[203] ^ x[89];
  assign t[163] = t[204] ^ x[90];
  assign t[164] = t[205] ^ x[91];
  assign t[165] = t[206] ^ x[92];
  assign t[166] = t[207] ^ x[93];
  assign t[167] = t[208] ^ x[94];
  assign t[168] = t[209] ^ x[95];
  assign t[169] = t[210] ^ x[96];
  assign t[16] = ~(t[103] & t[104]);
  assign t[170] = t[211] ^ x[97];
  assign t[171] = t[212] ^ x[98];
  assign t[172] = t[213] ^ x[104];
  assign t[173] = t[214] ^ x[105];
  assign t[174] = t[215] ^ x[106];
  assign t[175] = t[216] ^ x[107];
  assign t[176] = t[217] ^ x[108];
  assign t[177] = t[218] ^ x[109];
  assign t[178] = t[219] ^ x[110];
  assign t[179] = t[220] ^ x[111];
  assign t[17] = ~(t[105] & t[106]);
  assign t[180] = t[221] ^ x[112];
  assign t[181] = t[222] ^ x[113];
  assign t[182] = t[223] ^ x[114];
  assign t[183] = t[224] ^ x[115];
  assign t[184] = (~t[225] & t[226]);
  assign t[185] = (~t[227] & t[228]);
  assign t[186] = (~t[229] & t[230]);
  assign t[187] = (~t[231] & t[232]);
  assign t[188] = (~t[233] & t[234]);
  assign t[189] = (~t[235] & t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (~t[237] & t[238]);
  assign t[191] = (~t[235] & t[239]);
  assign t[192] = (~t[235] & t[240]);
  assign t[193] = (~t[241] & t[242]);
  assign t[194] = (~t[243] & t[244]);
  assign t[195] = (~t[237] & t[245]);
  assign t[196] = (~t[237] & t[246]);
  assign t[197] = (~t[247] & t[248]);
  assign t[198] = (~t[249] & t[250]);
  assign t[199] = (~t[251] & t[252]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[235] & t[253]);
  assign t[201] = (~t[241] & t[254]);
  assign t[202] = (~t[241] & t[255]);
  assign t[203] = (~t[256] & t[257]);
  assign t[204] = (~t[243] & t[258]);
  assign t[205] = (~t[243] & t[259]);
  assign t[206] = (~t[237] & t[260]);
  assign t[207] = (~t[247] & t[261]);
  assign t[208] = (~t[247] & t[262]);
  assign t[209] = (~t[249] & t[263]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[249] & t[264]);
  assign t[211] = (~t[251] & t[265]);
  assign t[212] = (~t[251] & t[266]);
  assign t[213] = (~t[267] & t[268]);
  assign t[214] = (~t[241] & t[269]);
  assign t[215] = (~t[256] & t[270]);
  assign t[216] = (~t[256] & t[271]);
  assign t[217] = (~t[243] & t[272]);
  assign t[218] = (~t[247] & t[273]);
  assign t[219] = (~t[249] & t[274]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[251] & t[275]);
  assign t[221] = (~t[267] & t[276]);
  assign t[222] = (~t[267] & t[277]);
  assign t[223] = (~t[256] & t[278]);
  assign t[224] = (~t[267] & t[279]);
  assign t[225] = t[280] ^ x[4];
  assign t[226] = t[281] ^ x[5];
  assign t[227] = t[282] ^ x[12];
  assign t[228] = t[283] ^ x[13];
  assign t[229] = t[284] ^ x[15];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[285] ^ x[16];
  assign t[231] = t[286] ^ x[18];
  assign t[232] = t[287] ^ x[19];
  assign t[233] = t[288] ^ x[21];
  assign t[234] = t[289] ^ x[22];
  assign t[235] = t[290] ^ x[27];
  assign t[236] = t[291] ^ x[28];
  assign t[237] = t[292] ^ x[35];
  assign t[238] = t[293] ^ x[36];
  assign t[239] = t[294] ^ x[39];
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = t[295] ^ x[40];
  assign t[241] = t[296] ^ x[45];
  assign t[242] = t[297] ^ x[46];
  assign t[243] = t[298] ^ x[53];
  assign t[244] = t[299] ^ x[54];
  assign t[245] = t[300] ^ x[57];
  assign t[246] = t[301] ^ x[58];
  assign t[247] = t[302] ^ x[63];
  assign t[248] = t[303] ^ x[64];
  assign t[249] = t[304] ^ x[69];
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = t[305] ^ x[70];
  assign t[251] = t[306] ^ x[77];
  assign t[252] = t[307] ^ x[78];
  assign t[253] = t[308] ^ x[81];
  assign t[254] = t[309] ^ x[82];
  assign t[255] = t[310] ^ x[83];
  assign t[256] = t[311] ^ x[88];
  assign t[257] = t[312] ^ x[89];
  assign t[258] = t[313] ^ x[90];
  assign t[259] = t[314] ^ x[91];
  assign t[25] = ~(t[105]);
  assign t[260] = t[315] ^ x[92];
  assign t[261] = t[316] ^ x[93];
  assign t[262] = t[317] ^ x[94];
  assign t[263] = t[318] ^ x[95];
  assign t[264] = t[319] ^ x[96];
  assign t[265] = t[320] ^ x[97];
  assign t[266] = t[321] ^ x[98];
  assign t[267] = t[322] ^ x[103];
  assign t[268] = t[323] ^ x[104];
  assign t[269] = t[324] ^ x[105];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[325] ^ x[106];
  assign t[271] = t[326] ^ x[107];
  assign t[272] = t[327] ^ x[108];
  assign t[273] = t[328] ^ x[109];
  assign t[274] = t[329] ^ x[110];
  assign t[275] = t[330] ^ x[111];
  assign t[276] = t[331] ^ x[112];
  assign t[277] = t[332] ^ x[113];
  assign t[278] = t[333] ^ x[114];
  assign t[279] = t[334] ^ x[115];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[281] = (x[3]);
  assign t[282] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[283] = (x[11]);
  assign t[284] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[285] = (x[14]);
  assign t[286] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[287] = (x[17]);
  assign t[288] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[289] = (x[20]);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[290] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[291] = (x[24]);
  assign t[292] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[293] = (x[32]);
  assign t[294] = (x[26]);
  assign t[295] = (x[23]);
  assign t[296] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[297] = (x[42]);
  assign t[298] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[299] = (x[50]);
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[34]);
  assign t[301] = (x[31]);
  assign t[302] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[303] = (x[60]);
  assign t[304] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[305] = (x[66]);
  assign t[306] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[307] = (x[74]);
  assign t[308] = (x[25]);
  assign t[309] = (x[44]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[41]);
  assign t[311] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[312] = (x[85]);
  assign t[313] = (x[52]);
  assign t[314] = (x[49]);
  assign t[315] = (x[33]);
  assign t[316] = (x[62]);
  assign t[317] = (x[59]);
  assign t[318] = (x[68]);
  assign t[319] = (x[65]);
  assign t[31] = t[47] | t[107];
  assign t[320] = (x[76]);
  assign t[321] = (x[73]);
  assign t[322] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[323] = (x[100]);
  assign t[324] = (x[43]);
  assign t[325] = (x[87]);
  assign t[326] = (x[84]);
  assign t[327] = (x[51]);
  assign t[328] = (x[61]);
  assign t[329] = (x[67]);
  assign t[32] = t[105] ? x[30] : x[29];
  assign t[330] = (x[75]);
  assign t[331] = (x[102]);
  assign t[332] = (x[99]);
  assign t[333] = (x[86]);
  assign t[334] = (x[101]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] ^ t[51];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[41];
  assign t[37] = ~(t[55] & t[56]);
  assign t[38] = t[57] | t[108];
  assign t[39] = t[18] ? x[38] : x[37];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[43];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[66];
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[110]);
  assign t[47] = ~(t[67] | t[45]);
  assign t[48] = ~(t[68] & t[69]);
  assign t[49] = t[70] | t[111];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[105] ? x[48] : x[47];
  assign t[51] = ~(t[71] & t[72]);
  assign t[52] = ~(t[73] & t[74]);
  assign t[53] = t[75] | t[112];
  assign t[54] = t[76] ? x[56] : x[55];
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[77] | t[55]);
  assign t[58] = ~(t[78] & t[79]);
  assign t[59] = t[80] | t[115];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[81] & t[82]);
  assign t[61] = t[83] | t[116];
  assign t[62] = t[76] ? x[72] : x[71];
  assign t[63] = ~(t[84] & t[85]);
  assign t[64] = t[86] | t[117];
  assign t[65] = t[76] ? x[80] : x[79];
  assign t[66] = ~(t[87] & t[88]);
  assign t[67] = ~(t[118]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[89] | t[68]);
  assign t[71] = ~(t[90] & t[91]);
  assign t[72] = t[92] | t[121];
  assign t[73] = ~(t[122]);
  assign t[74] = ~(t[123]);
  assign t[75] = ~(t[93] | t[73]);
  assign t[76] = ~(t[25]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[94] | t[78]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[95] | t[81]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[96] | t[84]);
  assign t[87] = ~(t[97] & t[98]);
  assign t[88] = t[99] | t[131];
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[100] | t[90]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[101] | t[97]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [115:0] x;
 output y;

 wire [343:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[139] & t[138]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[109] & t[110]);
  assign t[107] = ~(t[143] & t[142]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[5];
  assign t[153] = t[194] ^ x[13];
  assign t[154] = t[195] ^ x[16];
  assign t[155] = t[196] ^ x[19];
  assign t[156] = t[197] ^ x[22];
  assign t[157] = t[198] ^ x[28];
  assign t[158] = t[199] ^ x[36];
  assign t[159] = t[200] ^ x[39];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[40];
  assign t[161] = t[202] ^ x[46];
  assign t[162] = t[203] ^ x[54];
  assign t[163] = t[204] ^ x[57];
  assign t[164] = t[205] ^ x[58];
  assign t[165] = t[206] ^ x[64];
  assign t[166] = t[207] ^ x[70];
  assign t[167] = t[208] ^ x[78];
  assign t[168] = t[209] ^ x[81];
  assign t[169] = t[210] ^ x[82];
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = t[211] ^ x[83];
  assign t[171] = t[212] ^ x[89];
  assign t[172] = t[213] ^ x[90];
  assign t[173] = t[214] ^ x[91];
  assign t[174] = t[215] ^ x[92];
  assign t[175] = t[216] ^ x[93];
  assign t[176] = t[217] ^ x[94];
  assign t[177] = t[218] ^ x[95];
  assign t[178] = t[219] ^ x[96];
  assign t[179] = t[220] ^ x[97];
  assign t[17] = ~(t[114] & t[115]);
  assign t[180] = t[221] ^ x[98];
  assign t[181] = t[222] ^ x[104];
  assign t[182] = t[223] ^ x[105];
  assign t[183] = t[224] ^ x[106];
  assign t[184] = t[225] ^ x[107];
  assign t[185] = t[226] ^ x[108];
  assign t[186] = t[227] ^ x[109];
  assign t[187] = t[228] ^ x[110];
  assign t[188] = t[229] ^ x[111];
  assign t[189] = t[230] ^ x[112];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[113];
  assign t[191] = t[232] ^ x[114];
  assign t[192] = t[233] ^ x[115];
  assign t[193] = (~t[234] & t[235]);
  assign t[194] = (~t[236] & t[237]);
  assign t[195] = (~t[238] & t[239]);
  assign t[196] = (~t[240] & t[241]);
  assign t[197] = (~t[242] & t[243]);
  assign t[198] = (~t[244] & t[245]);
  assign t[199] = (~t[246] & t[247]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[244] & t[248]);
  assign t[201] = (~t[244] & t[249]);
  assign t[202] = (~t[250] & t[251]);
  assign t[203] = (~t[252] & t[253]);
  assign t[204] = (~t[246] & t[254]);
  assign t[205] = (~t[246] & t[255]);
  assign t[206] = (~t[256] & t[257]);
  assign t[207] = (~t[258] & t[259]);
  assign t[208] = (~t[260] & t[261]);
  assign t[209] = (~t[244] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[250] & t[263]);
  assign t[211] = (~t[250] & t[264]);
  assign t[212] = (~t[265] & t[266]);
  assign t[213] = (~t[252] & t[267]);
  assign t[214] = (~t[252] & t[268]);
  assign t[215] = (~t[246] & t[269]);
  assign t[216] = (~t[256] & t[270]);
  assign t[217] = (~t[256] & t[271]);
  assign t[218] = (~t[258] & t[272]);
  assign t[219] = (~t[258] & t[273]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[260] & t[274]);
  assign t[221] = (~t[260] & t[275]);
  assign t[222] = (~t[276] & t[277]);
  assign t[223] = (~t[250] & t[278]);
  assign t[224] = (~t[265] & t[279]);
  assign t[225] = (~t[265] & t[280]);
  assign t[226] = (~t[252] & t[281]);
  assign t[227] = (~t[256] & t[282]);
  assign t[228] = (~t[258] & t[283]);
  assign t[229] = (~t[260] & t[284]);
  assign t[22] = t[32] ^ t[21];
  assign t[230] = (~t[276] & t[285]);
  assign t[231] = (~t[276] & t[286]);
  assign t[232] = (~t[265] & t[287]);
  assign t[233] = (~t[276] & t[288]);
  assign t[234] = t[289] ^ x[4];
  assign t[235] = t[290] ^ x[5];
  assign t[236] = t[291] ^ x[12];
  assign t[237] = t[292] ^ x[13];
  assign t[238] = t[293] ^ x[15];
  assign t[239] = t[294] ^ x[16];
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = t[295] ^ x[18];
  assign t[241] = t[296] ^ x[19];
  assign t[242] = t[297] ^ x[21];
  assign t[243] = t[298] ^ x[22];
  assign t[244] = t[299] ^ x[27];
  assign t[245] = t[300] ^ x[28];
  assign t[246] = t[301] ^ x[35];
  assign t[247] = t[302] ^ x[36];
  assign t[248] = t[303] ^ x[39];
  assign t[249] = t[304] ^ x[40];
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = t[305] ^ x[45];
  assign t[251] = t[306] ^ x[46];
  assign t[252] = t[307] ^ x[53];
  assign t[253] = t[308] ^ x[54];
  assign t[254] = t[309] ^ x[57];
  assign t[255] = t[310] ^ x[58];
  assign t[256] = t[311] ^ x[63];
  assign t[257] = t[312] ^ x[64];
  assign t[258] = t[313] ^ x[69];
  assign t[259] = t[314] ^ x[70];
  assign t[25] = ~(t[114]);
  assign t[260] = t[315] ^ x[77];
  assign t[261] = t[316] ^ x[78];
  assign t[262] = t[317] ^ x[81];
  assign t[263] = t[318] ^ x[82];
  assign t[264] = t[319] ^ x[83];
  assign t[265] = t[320] ^ x[88];
  assign t[266] = t[321] ^ x[89];
  assign t[267] = t[322] ^ x[90];
  assign t[268] = t[323] ^ x[91];
  assign t[269] = t[324] ^ x[92];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[325] ^ x[93];
  assign t[271] = t[326] ^ x[94];
  assign t[272] = t[327] ^ x[95];
  assign t[273] = t[328] ^ x[96];
  assign t[274] = t[329] ^ x[97];
  assign t[275] = t[330] ^ x[98];
  assign t[276] = t[331] ^ x[103];
  assign t[277] = t[332] ^ x[104];
  assign t[278] = t[333] ^ x[105];
  assign t[279] = t[334] ^ x[106];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[335] ^ x[107];
  assign t[281] = t[336] ^ x[108];
  assign t[282] = t[337] ^ x[109];
  assign t[283] = t[338] ^ x[110];
  assign t[284] = t[339] ^ x[111];
  assign t[285] = t[340] ^ x[112];
  assign t[286] = t[341] ^ x[113];
  assign t[287] = t[342] ^ x[114];
  assign t[288] = t[343] ^ x[115];
  assign t[289] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[290] = (x[2]);
  assign t[291] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[292] = (x[11]);
  assign t[293] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[294] = (x[14]);
  assign t[295] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[296] = (x[17]);
  assign t[297] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[298] = (x[20]);
  assign t[299] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[24]);
  assign t[301] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[302] = (x[32]);
  assign t[303] = (x[26]);
  assign t[304] = (x[23]);
  assign t[305] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[306] = (x[42]);
  assign t[307] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[308] = (x[50]);
  assign t[309] = (x[34]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[31]);
  assign t[311] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[312] = (x[60]);
  assign t[313] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[314] = (x[66]);
  assign t[315] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[316] = (x[74]);
  assign t[317] = (x[25]);
  assign t[318] = (x[44]);
  assign t[319] = (x[41]);
  assign t[31] = ~(t[47] & t[116]);
  assign t[320] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[321] = (x[85]);
  assign t[322] = (x[52]);
  assign t[323] = (x[49]);
  assign t[324] = (x[33]);
  assign t[325] = (x[62]);
  assign t[326] = (x[59]);
  assign t[327] = (x[68]);
  assign t[328] = (x[65]);
  assign t[329] = (x[76]);
  assign t[32] = t[114] ? x[30] : x[29];
  assign t[330] = (x[73]);
  assign t[331] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[332] = (x[100]);
  assign t[333] = (x[43]);
  assign t[334] = (x[87]);
  assign t[335] = (x[84]);
  assign t[336] = (x[51]);
  assign t[337] = (x[61]);
  assign t[338] = (x[67]);
  assign t[339] = (x[75]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[102]);
  assign t[341] = (x[99]);
  assign t[342] = (x[86]);
  assign t[343] = (x[101]);
  assign t[34] = t[50] ^ t[51];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[41];
  assign t[37] = ~(t[55] & t[56]);
  assign t[38] = ~(t[57] & t[117]);
  assign t[39] = t[18] ? x[38] : x[37];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[43];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[66];
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[119]);
  assign t[47] = ~(t[67] & t[68]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = ~(t[71] & t[120]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[114] ? x[48] : x[47];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = ~(t[76] & t[121]);
  assign t[54] = t[18] ? x[56] : x[55];
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[77] & t[78]);
  assign t[58] = ~(t[79] & t[80]);
  assign t[59] = ~(t[81] & t[124]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = ~(t[84] & t[125]);
  assign t[62] = t[85] ? x[72] : x[71];
  assign t[63] = ~(t[86] & t[87]);
  assign t[64] = ~(t[88] & t[126]);
  assign t[65] = t[85] ? x[80] : x[79];
  assign t[66] = ~(t[89] & t[90]);
  assign t[67] = ~(t[119] & t[118]);
  assign t[68] = ~(t[127]);
  assign t[69] = ~(t[128]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[129]);
  assign t[71] = ~(t[91] & t[92]);
  assign t[72] = ~(t[93] & t[94]);
  assign t[73] = ~(t[95] & t[130]);
  assign t[74] = ~(t[131]);
  assign t[75] = ~(t[132]);
  assign t[76] = ~(t[96] & t[97]);
  assign t[77] = ~(t[123] & t[122]);
  assign t[78] = ~(t[133]);
  assign t[79] = ~(t[134]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[135]);
  assign t[81] = ~(t[98] & t[99]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[137]);
  assign t[84] = ~(t[100] & t[101]);
  assign t[85] = ~(t[25]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[102] & t[103]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[106] & t[140]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[143]);
  assign t[95] = ~(t[107] & t[108]);
  assign t[96] = ~(t[132] & t[131]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [106:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[5];
  assign t[127] = t[159] ^ x[13];
  assign t[128] = t[160] ^ x[16];
  assign t[129] = t[161] ^ x[19];
  assign t[12] = t[18] ? x[9] : x[10];
  assign t[130] = t[162] ^ x[22];
  assign t[131] = t[163] ^ x[28];
  assign t[132] = t[164] ^ x[29];
  assign t[133] = t[165] ^ x[37];
  assign t[134] = t[166] ^ x[38];
  assign t[135] = t[167] ^ x[41];
  assign t[136] = t[168] ^ x[47];
  assign t[137] = t[169] ^ x[48];
  assign t[138] = t[170] ^ x[56];
  assign t[139] = t[171] ^ x[57];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[60];
  assign t[141] = t[173] ^ x[66];
  assign t[142] = t[174] ^ x[67];
  assign t[143] = t[175] ^ x[73];
  assign t[144] = t[176] ^ x[74];
  assign t[145] = t[177] ^ x[82];
  assign t[146] = t[178] ^ x[83];
  assign t[147] = t[179] ^ x[86];
  assign t[148] = t[180] ^ x[92];
  assign t[149] = t[181] ^ x[93];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[94];
  assign t[151] = t[183] ^ x[95];
  assign t[152] = t[184] ^ x[96];
  assign t[153] = t[185] ^ x[102];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[104];
  assign t[156] = t[188] ^ x[105];
  assign t[157] = t[189] ^ x[106];
  assign t[158] = (~t[190] & t[191]);
  assign t[159] = (~t[192] & t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (~t[194] & t[195]);
  assign t[161] = (~t[196] & t[197]);
  assign t[162] = (~t[198] & t[199]);
  assign t[163] = (~t[200] & t[201]);
  assign t[164] = (~t[200] & t[202]);
  assign t[165] = (~t[203] & t[204]);
  assign t[166] = (~t[203] & t[205]);
  assign t[167] = (~t[200] & t[206]);
  assign t[168] = (~t[207] & t[208]);
  assign t[169] = (~t[207] & t[209]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (~t[210] & t[211]);
  assign t[171] = (~t[210] & t[212]);
  assign t[172] = (~t[203] & t[213]);
  assign t[173] = (~t[214] & t[215]);
  assign t[174] = (~t[214] & t[216]);
  assign t[175] = (~t[217] & t[218]);
  assign t[176] = (~t[217] & t[219]);
  assign t[177] = (~t[220] & t[221]);
  assign t[178] = (~t[220] & t[222]);
  assign t[179] = (~t[207] & t[223]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (~t[224] & t[225]);
  assign t[181] = (~t[224] & t[226]);
  assign t[182] = (~t[210] & t[227]);
  assign t[183] = (~t[214] & t[228]);
  assign t[184] = (~t[217] & t[229]);
  assign t[185] = (~t[230] & t[231]);
  assign t[186] = (~t[230] & t[232]);
  assign t[187] = (~t[220] & t[233]);
  assign t[188] = (~t[224] & t[234]);
  assign t[189] = (~t[230] & t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[236] ^ x[4];
  assign t[191] = t[237] ^ x[5];
  assign t[192] = t[238] ^ x[12];
  assign t[193] = t[239] ^ x[13];
  assign t[194] = t[240] ^ x[15];
  assign t[195] = t[241] ^ x[16];
  assign t[196] = t[242] ^ x[18];
  assign t[197] = t[243] ^ x[19];
  assign t[198] = t[244] ^ x[21];
  assign t[199] = t[245] ^ x[22];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[246] ^ x[27];
  assign t[201] = t[247] ^ x[28];
  assign t[202] = t[248] ^ x[29];
  assign t[203] = t[249] ^ x[36];
  assign t[204] = t[250] ^ x[37];
  assign t[205] = t[251] ^ x[38];
  assign t[206] = t[252] ^ x[41];
  assign t[207] = t[253] ^ x[46];
  assign t[208] = t[254] ^ x[47];
  assign t[209] = t[255] ^ x[48];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[256] ^ x[55];
  assign t[211] = t[257] ^ x[56];
  assign t[212] = t[258] ^ x[57];
  assign t[213] = t[259] ^ x[60];
  assign t[214] = t[260] ^ x[65];
  assign t[215] = t[261] ^ x[66];
  assign t[216] = t[262] ^ x[67];
  assign t[217] = t[263] ^ x[72];
  assign t[218] = t[264] ^ x[73];
  assign t[219] = t[265] ^ x[74];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[266] ^ x[81];
  assign t[221] = t[267] ^ x[82];
  assign t[222] = t[268] ^ x[83];
  assign t[223] = t[269] ^ x[86];
  assign t[224] = t[270] ^ x[91];
  assign t[225] = t[271] ^ x[92];
  assign t[226] = t[272] ^ x[93];
  assign t[227] = t[273] ^ x[94];
  assign t[228] = t[274] ^ x[95];
  assign t[229] = t[275] ^ x[96];
  assign t[22] = t[32] ^ t[21];
  assign t[230] = t[276] ^ x[101];
  assign t[231] = t[277] ^ x[102];
  assign t[232] = t[278] ^ x[103];
  assign t[233] = t[279] ^ x[104];
  assign t[234] = t[280] ^ x[105];
  assign t[235] = t[281] ^ x[106];
  assign t[236] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[237] = (x[1]);
  assign t[238] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[239] = (x[11]);
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[241] = (x[14]);
  assign t[242] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[243] = (x[17]);
  assign t[244] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[245] = (x[20]);
  assign t[246] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[247] = (x[25]);
  assign t[248] = (x[23]);
  assign t[249] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = (x[34]);
  assign t[251] = (x[32]);
  assign t[252] = (x[26]);
  assign t[253] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[254] = (x[44]);
  assign t[255] = (x[42]);
  assign t[256] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[257] = (x[53]);
  assign t[258] = (x[51]);
  assign t[259] = (x[35]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[261] = (x[63]);
  assign t[262] = (x[61]);
  assign t[263] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[264] = (x[70]);
  assign t[265] = (x[68]);
  assign t[266] = (x[77] & ~x[78] & ~x[79] & ~x[80]) | (~x[77] & x[78] & ~x[79] & ~x[80]) | (~x[77] & ~x[78] & x[79] & ~x[80]) | (~x[77] & ~x[78] & ~x[79] & x[80]) | (x[77] & x[78] & x[79] & ~x[80]) | (x[77] & x[78] & ~x[79] & x[80]) | (x[77] & ~x[78] & x[79] & x[80]) | (~x[77] & x[78] & x[79] & x[80]);
  assign t[267] = (x[79]);
  assign t[268] = (x[77]);
  assign t[269] = (x[45]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[87] & ~x[88] & ~x[89] & ~x[90]) | (~x[87] & x[88] & ~x[89] & ~x[90]) | (~x[87] & ~x[88] & x[89] & ~x[90]) | (~x[87] & ~x[88] & ~x[89] & x[90]) | (x[87] & x[88] & x[89] & ~x[90]) | (x[87] & x[88] & ~x[89] & x[90]) | (x[87] & ~x[88] & x[89] & x[90]) | (~x[87] & x[88] & x[89] & x[90]);
  assign t[271] = (x[89]);
  assign t[272] = (x[87]);
  assign t[273] = (x[54]);
  assign t[274] = (x[64]);
  assign t[275] = (x[71]);
  assign t[276] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[277] = (x[99]);
  assign t[278] = (x[97]);
  assign t[279] = (x[80]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[90]);
  assign t[281] = (x[100]);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[97] ? x[31] : x[30];
  assign t[33] = ~(t[47] & t[48]);
  assign t[34] = t[49] ^ t[50];
  assign t[35] = ~(t[51] & t[52]);
  assign t[36] = t[53] ^ t[43];
  assign t[37] = ~(t[101] & t[54]);
  assign t[38] = ~(t[102] & t[55]);
  assign t[39] = t[18] ? x[40] : x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[56] & t[57]);
  assign t[41] = ~(t[58] & t[59]);
  assign t[42] = t[60] ^ t[61];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[41];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[65]);
  assign t[47] = ~(t[104] & t[66]);
  assign t[48] = ~(t[105] & t[67]);
  assign t[49] = t[97] ? x[50] : x[49];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[68] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = ~(t[107] & t[71]);
  assign t[53] = t[72] ? x[59] : x[58];
  assign t[54] = ~(t[108]);
  assign t[55] = ~(t[108] & t[73]);
  assign t[56] = ~(t[109] & t[74]);
  assign t[57] = ~(t[110] & t[75]);
  assign t[58] = ~(t[111] & t[76]);
  assign t[59] = ~(t[112] & t[77]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[78] ? x[76] : x[75];
  assign t[61] = ~(t[79] & t[80]);
  assign t[62] = ~(t[113] & t[81]);
  assign t[63] = ~(t[114] & t[82]);
  assign t[64] = t[78] ? x[85] : x[84];
  assign t[65] = ~(t[99]);
  assign t[66] = ~(t[115]);
  assign t[67] = ~(t[115] & t[83]);
  assign t[68] = ~(t[116] & t[84]);
  assign t[69] = ~(t[117] & t[85]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[118]);
  assign t[71] = ~(t[118] & t[86]);
  assign t[72] = ~(t[25]);
  assign t[73] = ~(t[101]);
  assign t[74] = ~(t[119]);
  assign t[75] = ~(t[119] & t[87]);
  assign t[76] = ~(t[120]);
  assign t[77] = ~(t[120] & t[88]);
  assign t[78] = ~(t[25]);
  assign t[79] = ~(t[121] & t[89]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[122] & t[90]);
  assign t[81] = ~(t[123]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[124]);
  assign t[85] = ~(t[124] & t[92]);
  assign t[86] = ~(t[106]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[125]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125] & t[93]);
  assign t[91] = ~(t[113]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[121]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [115:0] x;
 output y;

 wire [427:0] t;
  assign t[0] = t[1] ? t[2] : t[195];
  assign t[100] = ~(t[217]);
  assign t[101] = ~(t[206] | t[207]);
  assign t[102] = ~(t[218]);
  assign t[103] = ~(t[219]);
  assign t[104] = ~(t[138] | t[139]);
  assign t[105] = ~(t[86] | t[140]);
  assign t[106] = ~(t[141] & t[142]);
  assign t[107] = ~(t[220]);
  assign t[108] = ~(t[221]);
  assign t[109] = ~(t[143] | t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[145] ? x[94] : x[93];
  assign t[111] = t[146] | t[147];
  assign t[112] = ~(t[222]);
  assign t[113] = ~(t[223]);
  assign t[114] = ~(t[148] | t[149]);
  assign t[115] = ~(t[150] | t[151]);
  assign t[116] = ~(t[224] | t[152]);
  assign t[117] = t[145] ? x[104] : x[103];
  assign t[118] = ~(t[153] & t[154]);
  assign t[119] = ~(t[198]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[155] & t[83]);
  assign t[121] = ~(t[156] & t[199]);
  assign t[122] = ~(t[119] | t[157]);
  assign t[123] = ~(t[79] | t[158]);
  assign t[124] = ~(t[159] & t[160]);
  assign t[125] = ~(t[161] & t[162]);
  assign t[126] = ~(t[163] | t[164]);
  assign t[127] = ~(t[165] | t[166]);
  assign t[128] = ~(t[225]);
  assign t[129] = ~(t[212] | t[213]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[163] | t[167]);
  assign t[131] = ~(t[168] | t[169]);
  assign t[132] = ~(t[226]);
  assign t[133] = ~(t[214] | t[215]);
  assign t[134] = ~(t[227]);
  assign t[135] = ~(t[228]);
  assign t[136] = ~(t[170] | t[171]);
  assign t[137] = ~(t[172] | t[166]);
  assign t[138] = ~(t[229]);
  assign t[139] = ~(t[218] | t[219]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = t[147] | t[164];
  assign t[141] = t[199] & t[161];
  assign t[142] = t[155] | t[156];
  assign t[143] = ~(t[230]);
  assign t[144] = ~(t[220] | t[221]);
  assign t[145] = ~(t[48]);
  assign t[146] = ~(t[173] & t[32]);
  assign t[147] = ~(t[79] | t[174]);
  assign t[148] = ~(t[231]);
  assign t[149] = ~(t[222] | t[223]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[232]);
  assign t[151] = ~(t[233]);
  assign t[152] = ~(t[175] | t[176]);
  assign t[153] = ~(t[49]);
  assign t[154] = ~(t[177] | t[147]);
  assign t[155] = ~(x[7] | t[197]);
  assign t[156] = x[7] & t[197];
  assign t[157] = t[196] ? t[120] : t[178];
  assign t[158] = t[196] ? t[180] : t[179];
  assign t[159] = ~(x[7] & t[181]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[199] & t[182]);
  assign t[161] = ~(t[119] | t[196]);
  assign t[162] = ~(t[160] & t[179]);
  assign t[163] = ~(t[79] | t[183]);
  assign t[164] = ~(t[79] | t[184]);
  assign t[165] = ~(t[79] | t[185]);
  assign t[166] = ~(t[79] | t[186]);
  assign t[167] = ~(t[187] & t[106]);
  assign t[168] = ~(t[119] | t[188]);
  assign t[169] = t[164] | t[189];
  assign t[16] = ~(t[196] & t[197]);
  assign t[170] = ~(t[234]);
  assign t[171] = ~(t[227] | t[228]);
  assign t[172] = ~(t[79] | t[190]);
  assign t[173] = ~(t[191] | t[168]);
  assign t[174] = t[196] ? t[160] : t[159];
  assign t[175] = ~(t[235]);
  assign t[176] = ~(t[232] | t[233]);
  assign t[177] = ~(t[137]);
  assign t[178] = ~(t[156] & t[83]);
  assign t[179] = ~(x[7] & t[51]);
  assign t[17] = ~(t[198] & t[199]);
  assign t[180] = ~(t[182] & t[83]);
  assign t[181] = ~(t[197] | t[199]);
  assign t[182] = ~(x[7] | t[192]);
  assign t[183] = t[196] ? t[120] : t[121];
  assign t[184] = t[196] ? t[193] : t[178];
  assign t[185] = t[196] ? t[159] : t[160];
  assign t[186] = t[196] ? t[178] : t[193];
  assign t[187] = ~(t[49] | t[165]);
  assign t[188] = t[196] ? t[180] : t[159];
  assign t[189] = ~(t[125]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = t[196] ? t[179] : t[180];
  assign t[191] = ~(t[119] | t[194]);
  assign t[192] = ~(t[197]);
  assign t[193] = ~(t[155] & t[199]);
  assign t[194] = t[196] ? t[178] : t[120];
  assign t[195] = (t[236]);
  assign t[196] = (t[237]);
  assign t[197] = (t[238]);
  assign t[198] = (t[239]);
  assign t[199] = (t[240]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = (t[241]);
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[9] : x[10];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = t[277] ^ x[5];
  assign t[237] = t[278] ^ x[13];
  assign t[238] = t[279] ^ x[16];
  assign t[239] = t[280] ^ x[19];
  assign t[23] = ~(t[22] ^ t[35]);
  assign t[240] = t[281] ^ x[22];
  assign t[241] = t[282] ^ x[28];
  assign t[242] = t[283] ^ x[34];
  assign t[243] = t[284] ^ x[35];
  assign t[244] = t[285] ^ x[36];
  assign t[245] = t[286] ^ x[44];
  assign t[246] = t[287] ^ x[50];
  assign t[247] = t[288] ^ x[51];
  assign t[248] = t[289] ^ x[52];
  assign t[249] = t[290] ^ x[58];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[66];
  assign t[251] = t[292] ^ x[72];
  assign t[252] = t[293] ^ x[73];
  assign t[253] = t[294] ^ x[74];
  assign t[254] = t[295] ^ x[75];
  assign t[255] = t[296] ^ x[78];
  assign t[256] = t[297] ^ x[79];
  assign t[257] = t[298] ^ x[85];
  assign t[258] = t[299] ^ x[88];
  assign t[259] = t[300] ^ x[89];
  assign t[25] = x[7] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[90];
  assign t[261] = t[302] ^ x[91];
  assign t[262] = t[303] ^ x[92];
  assign t[263] = t[304] ^ x[95];
  assign t[264] = t[305] ^ x[96];
  assign t[265] = t[306] ^ x[102];
  assign t[266] = t[307] ^ x[105];
  assign t[267] = t[308] ^ x[106];
  assign t[268] = t[309] ^ x[107];
  assign t[269] = t[310] ^ x[108];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[109];
  assign t[271] = t[312] ^ x[110];
  assign t[272] = t[313] ^ x[111];
  assign t[273] = t[314] ^ x[112];
  assign t[274] = t[315] ^ x[113];
  assign t[275] = t[316] ^ x[114];
  assign t[276] = t[317] ^ x[115];
  assign t[277] = (~t[318] & t[319]);
  assign t[278] = (~t[320] & t[321]);
  assign t[279] = (~t[322] & t[323]);
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = (~t[324] & t[325]);
  assign t[281] = (~t[326] & t[327]);
  assign t[282] = (~t[328] & t[329]);
  assign t[283] = (~t[330] & t[331]);
  assign t[284] = (~t[328] & t[332]);
  assign t[285] = (~t[328] & t[333]);
  assign t[286] = (~t[334] & t[335]);
  assign t[287] = (~t[336] & t[337]);
  assign t[288] = (~t[330] & t[338]);
  assign t[289] = (~t[330] & t[339]);
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = (~t[340] & t[341]);
  assign t[291] = (~t[342] & t[343]);
  assign t[292] = (~t[344] & t[345]);
  assign t[293] = (~t[328] & t[346]);
  assign t[294] = (~t[334] & t[347]);
  assign t[295] = (~t[334] & t[348]);
  assign t[296] = (~t[336] & t[349]);
  assign t[297] = (~t[336] & t[350]);
  assign t[298] = (~t[351] & t[352]);
  assign t[299] = (~t[330] & t[353]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[340] & t[354]);
  assign t[301] = (~t[340] & t[355]);
  assign t[302] = (~t[342] & t[356]);
  assign t[303] = (~t[342] & t[357]);
  assign t[304] = (~t[344] & t[358]);
  assign t[305] = (~t[344] & t[359]);
  assign t[306] = (~t[360] & t[361]);
  assign t[307] = (~t[334] & t[362]);
  assign t[308] = (~t[336] & t[363]);
  assign t[309] = (~t[351] & t[364]);
  assign t[30] = ~(t[48]);
  assign t[310] = (~t[351] & t[365]);
  assign t[311] = (~t[340] & t[366]);
  assign t[312] = (~t[342] & t[367]);
  assign t[313] = (~t[344] & t[368]);
  assign t[314] = (~t[360] & t[369]);
  assign t[315] = (~t[360] & t[370]);
  assign t[316] = (~t[351] & t[371]);
  assign t[317] = (~t[360] & t[372]);
  assign t[318] = t[373] ^ x[4];
  assign t[319] = t[374] ^ x[5];
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = t[375] ^ x[12];
  assign t[321] = t[376] ^ x[13];
  assign t[322] = t[377] ^ x[15];
  assign t[323] = t[378] ^ x[16];
  assign t[324] = t[379] ^ x[18];
  assign t[325] = t[380] ^ x[19];
  assign t[326] = t[381] ^ x[21];
  assign t[327] = t[382] ^ x[22];
  assign t[328] = t[383] ^ x[27];
  assign t[329] = t[384] ^ x[28];
  assign t[32] = ~(t[51] & t[52]);
  assign t[330] = t[385] ^ x[33];
  assign t[331] = t[386] ^ x[34];
  assign t[332] = t[387] ^ x[35];
  assign t[333] = t[388] ^ x[36];
  assign t[334] = t[389] ^ x[43];
  assign t[335] = t[390] ^ x[44];
  assign t[336] = t[391] ^ x[49];
  assign t[337] = t[392] ^ x[50];
  assign t[338] = t[393] ^ x[51];
  assign t[339] = t[394] ^ x[52];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[395] ^ x[57];
  assign t[341] = t[396] ^ x[58];
  assign t[342] = t[397] ^ x[65];
  assign t[343] = t[398] ^ x[66];
  assign t[344] = t[399] ^ x[71];
  assign t[345] = t[400] ^ x[72];
  assign t[346] = t[401] ^ x[73];
  assign t[347] = t[402] ^ x[74];
  assign t[348] = t[403] ^ x[75];
  assign t[349] = t[404] ^ x[78];
  assign t[34] = ~(t[200] | t[55]);
  assign t[350] = t[405] ^ x[79];
  assign t[351] = t[406] ^ x[84];
  assign t[352] = t[407] ^ x[85];
  assign t[353] = t[408] ^ x[88];
  assign t[354] = t[409] ^ x[89];
  assign t[355] = t[410] ^ x[90];
  assign t[356] = t[411] ^ x[91];
  assign t[357] = t[412] ^ x[92];
  assign t[358] = t[413] ^ x[95];
  assign t[359] = t[414] ^ x[96];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[415] ^ x[101];
  assign t[361] = t[416] ^ x[102];
  assign t[362] = t[417] ^ x[105];
  assign t[363] = t[418] ^ x[106];
  assign t[364] = t[419] ^ x[107];
  assign t[365] = t[420] ^ x[108];
  assign t[366] = t[421] ^ x[109];
  assign t[367] = t[422] ^ x[110];
  assign t[368] = t[423] ^ x[111];
  assign t[369] = t[424] ^ x[112];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[425] ^ x[113];
  assign t[371] = t[426] ^ x[114];
  assign t[372] = t[427] ^ x[115];
  assign t[373] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[374] = (x[0]);
  assign t[375] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[376] = (x[11]);
  assign t[377] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[378] = (x[14]);
  assign t[379] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = ~(t[44] ^ t[60]);
  assign t[380] = (x[17]);
  assign t[381] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[382] = (x[20]);
  assign t[383] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[384] = (x[24]);
  assign t[385] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[386] = (x[30]);
  assign t[387] = (x[25]);
  assign t[388] = (x[26]);
  assign t[389] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[38] = ~(t[61] | t[62]);
  assign t[390] = (x[40]);
  assign t[391] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[392] = (x[46]);
  assign t[393] = (x[31]);
  assign t[394] = (x[32]);
  assign t[395] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[396] = (x[54]);
  assign t[397] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[398] = (x[62]);
  assign t[399] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[39] = ~(t[63] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[68]);
  assign t[401] = (x[23]);
  assign t[402] = (x[41]);
  assign t[403] = (x[42]);
  assign t[404] = (x[47]);
  assign t[405] = (x[48]);
  assign t[406] = (x[80] & ~x[81] & ~x[82] & ~x[83]) | (~x[80] & x[81] & ~x[82] & ~x[83]) | (~x[80] & ~x[81] & x[82] & ~x[83]) | (~x[80] & ~x[81] & ~x[82] & x[83]) | (x[80] & x[81] & x[82] & ~x[83]) | (x[80] & x[81] & ~x[82] & x[83]) | (x[80] & ~x[81] & x[82] & x[83]) | (~x[80] & x[81] & x[82] & x[83]);
  assign t[407] = (x[81]);
  assign t[408] = (x[29]);
  assign t[409] = (x[55]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[56]);
  assign t[411] = (x[63]);
  assign t[412] = (x[64]);
  assign t[413] = (x[69]);
  assign t[414] = (x[70]);
  assign t[415] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[416] = (x[98]);
  assign t[417] = (x[39]);
  assign t[418] = (x[45]);
  assign t[419] = (x[82]);
  assign t[41] = ~(t[201] | t[67]);
  assign t[420] = (x[83]);
  assign t[421] = (x[53]);
  assign t[422] = (x[61]);
  assign t[423] = (x[67]);
  assign t[424] = (x[99]);
  assign t[425] = (x[100]);
  assign t[426] = (x[80]);
  assign t[427] = (x[97]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[45] = ~(t[46] ^ t[74]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[48] = ~(t[198]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[81] & t[82]);
  assign t[51] = ~(t[197] | t[83]);
  assign t[52] = t[79] & t[196];
  assign t[53] = ~(t[202]);
  assign t[54] = ~(t[203]);
  assign t[55] = ~(t[84] | t[85]);
  assign t[56] = t[198] ? x[38] : x[37];
  assign t[57] = t[86] | t[87];
  assign t[58] = ~(t[88] | t[89]);
  assign t[59] = ~(t[204] | t[90]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[91] ^ t[92]);
  assign t[61] = ~(t[93] | t[94]);
  assign t[62] = ~(t[205] | t[95]);
  assign t[63] = ~(t[96] | t[97]);
  assign t[64] = ~(t[98] ^ t[99]);
  assign t[65] = ~(t[206]);
  assign t[66] = ~(t[207]);
  assign t[67] = ~(t[100] | t[101]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[208] | t[104]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[30] ? x[60] : x[59];
  assign t[71] = ~(t[105] & t[106]);
  assign t[72] = ~(t[107] | t[108]);
  assign t[73] = ~(t[209] | t[109]);
  assign t[74] = ~(t[110] ^ t[111]);
  assign t[75] = ~(t[112] | t[113]);
  assign t[76] = ~(t[210] | t[114]);
  assign t[77] = ~(t[115] | t[116]);
  assign t[78] = ~(t[117] ^ t[118]);
  assign t[79] = ~(t[119]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[196] ? t[121] : t[120];
  assign t[81] = ~(t[122] | t[123]);
  assign t[82] = ~(t[119] & t[124]);
  assign t[83] = ~(t[199]);
  assign t[84] = ~(t[211]);
  assign t[85] = ~(t[202] | t[203]);
  assign t[86] = ~(t[125] & t[32]);
  assign t[87] = ~(t[126] & t[127]);
  assign t[88] = ~(t[212]);
  assign t[89] = ~(t[213]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[128] | t[129]);
  assign t[91] = t[198] ? x[77] : x[76];
  assign t[92] = ~(t[130] & t[131]);
  assign t[93] = ~(t[214]);
  assign t[94] = ~(t[215]);
  assign t[95] = ~(t[132] | t[133]);
  assign t[96] = ~(t[134] | t[135]);
  assign t[97] = ~(t[216] | t[136]);
  assign t[98] = t[198] ? x[87] : x[86];
  assign t[99] = ~(t[130] & t[137]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [172:0] x;
 output y;

 wire [673:0] t;
  assign t[0] = t[1] ? t[2] : t[404];
  assign t[100] = ~(t[426] | t[142]);
  assign t[101] = t[30] ? x[91] : x[90];
  assign t[102] = ~(t[143] & t[144]);
  assign t[103] = ~(t[427]);
  assign t[104] = ~(t[428]);
  assign t[105] = ~(t[145] | t[146]);
  assign t[106] = t[30] ? x[95] : x[94];
  assign t[107] = ~(t[147] & t[148]);
  assign t[108] = ~(t[429]);
  assign t[109] = ~(t[416] | t[417]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[430]);
  assign t[111] = ~(t[431]);
  assign t[112] = ~(t[149] | t[150]);
  assign t[113] = ~(t[151] | t[152]);
  assign t[114] = ~(t[432]);
  assign t[115] = ~(t[433]);
  assign t[116] = ~(t[153] | t[154]);
  assign t[117] = t[155] ? x[102] : x[101];
  assign t[118] = t[156] | t[84];
  assign t[119] = ~(t[434]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[435]);
  assign t[121] = ~(t[157] | t[158]);
  assign t[122] = ~(t[159] | t[160]);
  assign t[123] = ~(t[436] | t[161]);
  assign t[124] = t[155] ? x[112] : x[111];
  assign t[125] = ~(t[162] & t[163]);
  assign t[126] = ~(t[164] & t[165]);
  assign t[127] = ~(t[406] | t[166]);
  assign t[128] = t[129] & t[405];
  assign t[129] = ~(t[132]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[405] ? t[164] : t[167];
  assign t[131] = t[405] ? t[169] : t[168];
  assign t[132] = ~(t[407]);
  assign t[133] = ~(t[437]);
  assign t[134] = ~(t[422] | t[423]);
  assign t[135] = ~(t[132] | t[170]);
  assign t[136] = ~(t[129] | t[171]);
  assign t[137] = ~(t[172] & t[173]);
  assign t[138] = ~(t[438]);
  assign t[139] = ~(t[424] | t[425]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[439]);
  assign t[141] = ~(t[440]);
  assign t[142] = ~(t[174] | t[175]);
  assign t[143] = ~(t[151] | t[176]);
  assign t[144] = ~(t[118] | t[177]);
  assign t[145] = ~(t[441]);
  assign t[146] = ~(t[427] | t[428]);
  assign t[147] = ~(t[178] | t[85]);
  assign t[148] = ~(t[135] | t[156]);
  assign t[149] = ~(t[442]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[430] | t[431]);
  assign t[151] = ~(t[129] | t[179]);
  assign t[152] = ~(t[94] & t[180]);
  assign t[153] = ~(t[443]);
  assign t[154] = ~(t[432] | t[433]);
  assign t[155] = ~(t[49]);
  assign t[156] = ~(t[181] & t[83]);
  assign t[157] = ~(t[444]);
  assign t[158] = ~(t[434] | t[435]);
  assign t[159] = ~(t[445]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[446]);
  assign t[161] = ~(t[182] | t[183]);
  assign t[162] = ~(t[151]);
  assign t[163] = ~(t[184] | t[84]);
  assign t[164] = ~(t[408] & t[185]);
  assign t[165] = ~(x[7] & t[127]);
  assign t[166] = ~(t[408]);
  assign t[167] = ~(x[7] & t[186]);
  assign t[168] = ~(t[88] & t[166]);
  assign t[169] = ~(t[87] & t[408]);
  assign t[16] = ~(t[405] & t[406]);
  assign t[170] = t[405] ? t[187] : t[168];
  assign t[171] = t[405] ? t[188] : t[165];
  assign t[172] = ~(t[151] | t[189]);
  assign t[173] = t[132] | t[190];
  assign t[174] = ~(t[447]);
  assign t[175] = ~(t[439] | t[440]);
  assign t[176] = ~(t[129] | t[191]);
  assign t[177] = ~(t[192] & t[173]);
  assign t[178] = ~(t[129] | t[193]);
  assign t[179] = t[405] ? t[194] : t[187];
  assign t[17] = ~(t[407] & t[408]);
  assign t[180] = ~(t[132] & t[195]);
  assign t[181] = ~(t[196] | t[197]);
  assign t[182] = ~(t[448]);
  assign t[183] = ~(t[445] | t[446]);
  assign t[184] = ~(t[198]);
  assign t[185] = ~(x[7] | t[199]);
  assign t[186] = ~(t[406] | t[408]);
  assign t[187] = ~(t[87] & t[166]);
  assign t[188] = ~(t[185] & t[166]);
  assign t[189] = ~(t[129] | t[200]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = t[405] ? t[167] : t[188];
  assign t[191] = t[405] ? t[167] : t[164];
  assign t[192] = ~(t[201] | t[202]);
  assign t[193] = t[405] ? t[187] : t[194];
  assign t[194] = ~(t[88] & t[408]);
  assign t[195] = ~(t[167] & t[164]);
  assign t[196] = ~(t[132] | t[203]);
  assign t[197] = ~(t[132] | t[204]);
  assign t[198] = ~(t[202] | t[189]);
  assign t[199] = ~(t[406]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[405] ? t[168] : t[169];
  assign t[201] = ~(t[82]);
  assign t[202] = ~(t[129] | t[205]);
  assign t[203] = t[405] ? t[168] : t[187];
  assign t[204] = t[405] ? t[188] : t[167];
  assign t[205] = t[405] ? t[165] : t[188];
  assign t[206] = t[1] ? t[207] : t[449];
  assign t[207] = x[6] ? t[209] : t[208];
  assign t[208] = x[7] ? t[211] : t[210];
  assign t[209] = t[212] ^ x[126];
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = t[213] ^ t[214];
  assign t[211] = ~(t[215] ^ t[216]);
  assign t[212] = x[127] ^ x[128];
  assign t[213] = t[30] ? x[128] : x[127];
  assign t[214] = ~(t[217] ^ t[218]);
  assign t[215] = x[7] ? t[220] : t[219];
  assign t[216] = ~(t[221] ^ t[222]);
  assign t[217] = x[7] ? t[224] : t[223];
  assign t[218] = ~(t[225] ^ t[226]);
  assign t[219] = ~(t[227] & t[228]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = t[229] ^ t[230];
  assign t[221] = x[7] ? t[232] : t[231];
  assign t[222] = x[7] ? t[234] : t[233];
  assign t[223] = ~(t[235] & t[236]);
  assign t[224] = t[237] ^ t[238];
  assign t[225] = x[7] ? t[240] : t[239];
  assign t[226] = x[7] ? t[242] : t[241];
  assign t[227] = ~(t[411] & t[55]);
  assign t[228] = ~(t[421] & t[243]);
  assign t[229] = t[30] ? x[130] : x[129];
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = ~(t[244] & t[245]);
  assign t[231] = ~(t[246] & t[247]);
  assign t[232] = t[248] ^ t[233];
  assign t[233] = ~(t[249] & t[250]);
  assign t[234] = t[251] ^ t[252];
  assign t[235] = ~(t[416] & t[69]);
  assign t[236] = ~(t[429] & t[253]);
  assign t[237] = t[30] ? x[132] : x[131];
  assign t[238] = ~(t[254] & t[255]);
  assign t[239] = ~(t[256] & t[257]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = t[258] ^ t[259];
  assign t[241] = ~(t[260] & t[261]);
  assign t[242] = t[262] ^ t[239];
  assign t[243] = ~(t[412] & t[54]);
  assign t[244] = ~(t[422] & t[92]);
  assign t[245] = ~(t[437] & t[263]);
  assign t[246] = ~(t[427] & t[104]);
  assign t[247] = ~(t[441] & t[264]);
  assign t[248] = t[155] ? x[134] : x[133];
  assign t[249] = ~(t[424] & t[97]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = ~(t[438] & t[265]);
  assign t[251] = t[30] ? x[136] : x[135];
  assign t[252] = ~(t[266] & t[267]);
  assign t[253] = ~(t[417] & t[68]);
  assign t[254] = ~(t[430] & t[111]);
  assign t[255] = ~(t[442] & t[268]);
  assign t[256] = ~(t[434] & t[120]);
  assign t[257] = ~(t[444] & t[269]);
  assign t[258] = t[155] ? x[138] : x[137];
  assign t[259] = ~(t[270] & t[271]);
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = ~(t[432] & t[115]);
  assign t[261] = ~(t[443] & t[272]);
  assign t[262] = t[155] ? x[140] : x[139];
  assign t[263] = ~(t[423] & t[91]);
  assign t[264] = ~(t[428] & t[103]);
  assign t[265] = ~(t[425] & t[96]);
  assign t[266] = ~(t[439] & t[141]);
  assign t[267] = ~(t[447] & t[273]);
  assign t[268] = ~(t[431] & t[110]);
  assign t[269] = ~(t[435] & t[119]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = ~(t[445] & t[160]);
  assign t[271] = ~(t[448] & t[274]);
  assign t[272] = ~(t[433] & t[114]);
  assign t[273] = ~(t[440] & t[140]);
  assign t[274] = ~(t[446] & t[159]);
  assign t[275] = t[1] ? t[276] : t[450];
  assign t[276] = x[6] ? t[278] : t[277];
  assign t[277] = x[7] ? t[280] : t[279];
  assign t[278] = t[281] ^ x[142];
  assign t[279] = t[282] ^ t[283];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = ~(t[284] ^ t[285]);
  assign t[281] = x[143] ^ x[144];
  assign t[282] = t[30] ? x[144] : x[143];
  assign t[283] = ~(t[286] ^ t[287]);
  assign t[284] = x[7] ? t[289] : t[288];
  assign t[285] = ~(t[290] ^ t[291]);
  assign t[286] = x[7] ? t[293] : t[292];
  assign t[287] = ~(t[294] ^ t[295]);
  assign t[288] = ~(t[296] & t[297]);
  assign t[289] = t[298] ^ t[299];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = x[7] ? t[301] : t[300];
  assign t[291] = x[7] ? t[303] : t[302];
  assign t[292] = ~(t[304] & t[305]);
  assign t[293] = t[306] ^ t[307];
  assign t[294] = x[7] ? t[309] : t[308];
  assign t[295] = x[7] ? t[311] : t[310];
  assign t[296] = ~(t[55] & t[89]);
  assign t[297] = ~(t[312] & t[409]);
  assign t[298] = t[155] ? x[146] : x[145];
  assign t[299] = ~(t[313] & t[314]);
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = ~(t[315] & t[316]);
  assign t[301] = t[317] ^ t[318];
  assign t[302] = ~(t[319] & t[320]);
  assign t[303] = t[321] ^ t[300];
  assign t[304] = ~(t[69] & t[108]);
  assign t[305] = ~(t[322] & t[410]);
  assign t[306] = t[30] ? x[148] : x[147];
  assign t[307] = ~(t[323] & t[324]);
  assign t[308] = ~(t[325] & t[326]);
  assign t[309] = t[327] ^ t[310];
  assign t[30] = ~(t[49]);
  assign t[310] = ~(t[328] & t[329]);
  assign t[311] = t[330] ^ t[331];
  assign t[312] = ~(t[332] & t[54]);
  assign t[313] = ~(t[92] & t[133]);
  assign t[314] = ~(t[333] & t[413]);
  assign t[315] = ~(t[97] & t[138]);
  assign t[316] = ~(t[334] & t[414]);
  assign t[317] = t[30] ? x[150] : x[149];
  assign t[318] = ~(t[335] & t[336]);
  assign t[319] = ~(t[104] & t[145]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = ~(t[337] & t[415]);
  assign t[321] = t[407] ? x[152] : x[151];
  assign t[322] = ~(t[338] & t[68]);
  assign t[323] = ~(t[111] & t[149]);
  assign t[324] = ~(t[339] & t[418]);
  assign t[325] = ~(t[115] & t[153]);
  assign t[326] = ~(t[340] & t[419]);
  assign t[327] = t[155] ? x[154] : x[153];
  assign t[328] = ~(t[120] & t[157]);
  assign t[329] = ~(t[341] & t[420]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[330] = t[155] ? x[156] : x[155];
  assign t[331] = ~(t[342] & t[343]);
  assign t[332] = ~(t[421] & t[412]);
  assign t[333] = ~(t[344] & t[91]);
  assign t[334] = ~(t[345] & t[96]);
  assign t[335] = ~(t[141] & t[174]);
  assign t[336] = ~(t[346] & t[426]);
  assign t[337] = ~(t[347] & t[103]);
  assign t[338] = ~(t[429] & t[417]);
  assign t[339] = ~(t[348] & t[110]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = ~(t[349] & t[114]);
  assign t[341] = ~(t[350] & t[119]);
  assign t[342] = ~(t[160] & t[182]);
  assign t[343] = ~(t[351] & t[436]);
  assign t[344] = ~(t[437] & t[423]);
  assign t[345] = ~(t[438] & t[425]);
  assign t[346] = ~(t[352] & t[140]);
  assign t[347] = ~(t[441] & t[428]);
  assign t[348] = ~(t[442] & t[431]);
  assign t[349] = ~(t[443] & t[433]);
  assign t[34] = ~(t[409] | t[56]);
  assign t[350] = ~(t[444] & t[435]);
  assign t[351] = ~(t[353] & t[159]);
  assign t[352] = ~(t[447] & t[440]);
  assign t[353] = ~(t[448] & t[446]);
  assign t[354] = t[1] ? t[355] : t[451];
  assign t[355] = x[6] ? t[357] : t[356];
  assign t[356] = x[7] ? t[359] : t[358];
  assign t[357] = t[360] ^ x[158];
  assign t[358] = t[361] ^ t[362];
  assign t[359] = ~(t[363] ^ t[364]);
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = x[159] ^ x[160];
  assign t[361] = t[30] ? x[160] : x[159];
  assign t[362] = ~(t[365] ^ t[366]);
  assign t[363] = x[7] ? t[368] : t[367];
  assign t[364] = ~(t[369] ^ t[370]);
  assign t[365] = x[7] ? t[372] : t[371];
  assign t[366] = ~(t[373] ^ t[374]);
  assign t[367] = ~(t[296] & t[375]);
  assign t[368] = t[376] ^ t[377];
  assign t[369] = x[7] ? t[379] : t[378];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = x[7] ? t[381] : t[380];
  assign t[371] = ~(t[304] & t[382]);
  assign t[372] = t[383] ^ t[384];
  assign t[373] = x[7] ? t[386] : t[385];
  assign t[374] = x[7] ? t[388] : t[387];
  assign t[375] = t[33] | t[409];
  assign t[376] = t[389] ? x[162] : x[161];
  assign t[377] = ~(t[313] & t[390]);
  assign t[378] = ~(t[315] & t[391]);
  assign t[379] = t[392] ^ t[393];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = ~(t[319] & t[394]);
  assign t[381] = t[395] ^ t[378];
  assign t[382] = t[41] | t[410];
  assign t[383] = t[30] ? x[164] : x[163];
  assign t[384] = ~(t[323] & t[396]);
  assign t[385] = ~(t[325] & t[397]);
  assign t[386] = t[398] ^ t[387];
  assign t[387] = ~(t[328] & t[399]);
  assign t[388] = t[400] ^ t[401];
  assign t[389] = ~(t[49]);
  assign t[38] = ~(t[63] ^ t[64]);
  assign t[390] = t[57] | t[413];
  assign t[391] = t[61] | t[414];
  assign t[392] = t[30] ? x[166] : x[165];
  assign t[393] = ~(t[335] & t[402]);
  assign t[394] = t[65] | t[415];
  assign t[395] = t[30] ? x[168] : x[167];
  assign t[396] = t[71] | t[418];
  assign t[397] = t[75] | t[419];
  assign t[398] = t[155] ? x[170] : x[169];
  assign t[399] = t[78] | t[420];
  assign t[39] = ~(t[65] | t[66]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[155] ? x[172] : x[171];
  assign t[401] = ~(t[342] & t[403]);
  assign t[402] = t[99] | t[426];
  assign t[403] = t[122] | t[436];
  assign t[404] = (t[452]);
  assign t[405] = (t[453]);
  assign t[406] = (t[454]);
  assign t[407] = (t[455]);
  assign t[408] = (t[456]);
  assign t[409] = (t[457]);
  assign t[40] = ~(t[37] ^ t[67]);
  assign t[410] = (t[458]);
  assign t[411] = (t[459]);
  assign t[412] = (t[460]);
  assign t[413] = (t[461]);
  assign t[414] = (t[462]);
  assign t[415] = (t[463]);
  assign t[416] = (t[464]);
  assign t[417] = (t[465]);
  assign t[418] = (t[466]);
  assign t[419] = (t[467]);
  assign t[41] = ~(t[68] | t[69]);
  assign t[420] = (t[468]);
  assign t[421] = (t[469]);
  assign t[422] = (t[470]);
  assign t[423] = (t[471]);
  assign t[424] = (t[472]);
  assign t[425] = (t[473]);
  assign t[426] = (t[474]);
  assign t[427] = (t[475]);
  assign t[428] = (t[476]);
  assign t[429] = (t[477]);
  assign t[42] = ~(t[410] | t[70]);
  assign t[430] = (t[478]);
  assign t[431] = (t[479]);
  assign t[432] = (t[480]);
  assign t[433] = (t[481]);
  assign t[434] = (t[482]);
  assign t[435] = (t[483]);
  assign t[436] = (t[484]);
  assign t[437] = (t[485]);
  assign t[438] = (t[486]);
  assign t[439] = (t[487]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[440] = (t[488]);
  assign t[441] = (t[489]);
  assign t[442] = (t[490]);
  assign t[443] = (t[491]);
  assign t[444] = (t[492]);
  assign t[445] = (t[493]);
  assign t[446] = (t[494]);
  assign t[447] = (t[495]);
  assign t[448] = (t[496]);
  assign t[449] = (t[497]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[450] = (t[498]);
  assign t[451] = (t[499]);
  assign t[452] = t[500] ^ x[5];
  assign t[453] = t[501] ^ x[13];
  assign t[454] = t[502] ^ x[16];
  assign t[455] = t[503] ^ x[19];
  assign t[456] = t[504] ^ x[22];
  assign t[457] = t[505] ^ x[28];
  assign t[458] = t[506] ^ x[34];
  assign t[459] = t[507] ^ x[35];
  assign t[45] = ~(t[75] | t[76]);
  assign t[460] = t[508] ^ x[36];
  assign t[461] = t[509] ^ x[42];
  assign t[462] = t[510] ^ x[50];
  assign t[463] = t[511] ^ x[56];
  assign t[464] = t[512] ^ x[57];
  assign t[465] = t[513] ^ x[58];
  assign t[466] = t[514] ^ x[64];
  assign t[467] = t[515] ^ x[72];
  assign t[468] = t[516] ^ x[78];
  assign t[469] = t[517] ^ x[79];
  assign t[46] = ~(t[47] ^ t[77]);
  assign t[470] = t[518] ^ x[80];
  assign t[471] = t[519] ^ x[81];
  assign t[472] = t[520] ^ x[82];
  assign t[473] = t[521] ^ x[83];
  assign t[474] = t[522] ^ x[89];
  assign t[475] = t[523] ^ x[92];
  assign t[476] = t[524] ^ x[93];
  assign t[477] = t[525] ^ x[96];
  assign t[478] = t[526] ^ x[97];
  assign t[479] = t[527] ^ x[98];
  assign t[47] = ~(t[78] | t[79]);
  assign t[480] = t[528] ^ x[99];
  assign t[481] = t[529] ^ x[100];
  assign t[482] = t[530] ^ x[103];
  assign t[483] = t[531] ^ x[104];
  assign t[484] = t[532] ^ x[110];
  assign t[485] = t[533] ^ x[113];
  assign t[486] = t[534] ^ x[114];
  assign t[487] = t[535] ^ x[115];
  assign t[488] = t[536] ^ x[116];
  assign t[489] = t[537] ^ x[117];
  assign t[48] = ~(t[80] ^ t[81]);
  assign t[490] = t[538] ^ x[118];
  assign t[491] = t[539] ^ x[119];
  assign t[492] = t[540] ^ x[120];
  assign t[493] = t[541] ^ x[121];
  assign t[494] = t[542] ^ x[122];
  assign t[495] = t[543] ^ x[123];
  assign t[496] = t[544] ^ x[124];
  assign t[497] = t[545] ^ x[125];
  assign t[498] = t[546] ^ x[141];
  assign t[499] = t[547] ^ x[157];
  assign t[49] = ~(t[407]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[548] & t[549]);
  assign t[501] = (~t[550] & t[551]);
  assign t[502] = (~t[552] & t[553]);
  assign t[503] = (~t[554] & t[555]);
  assign t[504] = (~t[556] & t[557]);
  assign t[505] = (~t[558] & t[559]);
  assign t[506] = (~t[560] & t[561]);
  assign t[507] = (~t[558] & t[562]);
  assign t[508] = (~t[558] & t[563]);
  assign t[509] = (~t[564] & t[565]);
  assign t[50] = ~(t[82] & t[83]);
  assign t[510] = (~t[566] & t[567]);
  assign t[511] = (~t[568] & t[569]);
  assign t[512] = (~t[560] & t[570]);
  assign t[513] = (~t[560] & t[571]);
  assign t[514] = (~t[572] & t[573]);
  assign t[515] = (~t[574] & t[575]);
  assign t[516] = (~t[576] & t[577]);
  assign t[517] = (~t[558] & t[578]);
  assign t[518] = (~t[564] & t[579]);
  assign t[519] = (~t[564] & t[580]);
  assign t[51] = t[84] | t[85];
  assign t[520] = (~t[566] & t[581]);
  assign t[521] = (~t[566] & t[582]);
  assign t[522] = (~t[583] & t[584]);
  assign t[523] = (~t[568] & t[585]);
  assign t[524] = (~t[568] & t[586]);
  assign t[525] = (~t[560] & t[587]);
  assign t[526] = (~t[572] & t[588]);
  assign t[527] = (~t[572] & t[589]);
  assign t[528] = (~t[574] & t[590]);
  assign t[529] = (~t[574] & t[591]);
  assign t[52] = t[408] & t[86];
  assign t[530] = (~t[576] & t[592]);
  assign t[531] = (~t[576] & t[593]);
  assign t[532] = (~t[594] & t[595]);
  assign t[533] = (~t[564] & t[596]);
  assign t[534] = (~t[566] & t[597]);
  assign t[535] = (~t[583] & t[598]);
  assign t[536] = (~t[583] & t[599]);
  assign t[537] = (~t[568] & t[600]);
  assign t[538] = (~t[572] & t[601]);
  assign t[539] = (~t[574] & t[602]);
  assign t[53] = t[87] | t[88];
  assign t[540] = (~t[576] & t[603]);
  assign t[541] = (~t[594] & t[604]);
  assign t[542] = (~t[594] & t[605]);
  assign t[543] = (~t[583] & t[606]);
  assign t[544] = (~t[594] & t[607]);
  assign t[545] = (~t[548] & t[608]);
  assign t[546] = (~t[548] & t[609]);
  assign t[547] = (~t[548] & t[610]);
  assign t[548] = t[611] ^ x[4];
  assign t[549] = t[612] ^ x[5];
  assign t[54] = ~(t[411]);
  assign t[550] = t[613] ^ x[12];
  assign t[551] = t[614] ^ x[13];
  assign t[552] = t[615] ^ x[15];
  assign t[553] = t[616] ^ x[16];
  assign t[554] = t[617] ^ x[18];
  assign t[555] = t[618] ^ x[19];
  assign t[556] = t[619] ^ x[21];
  assign t[557] = t[620] ^ x[22];
  assign t[558] = t[621] ^ x[27];
  assign t[559] = t[622] ^ x[28];
  assign t[55] = ~(t[412]);
  assign t[560] = t[623] ^ x[33];
  assign t[561] = t[624] ^ x[34];
  assign t[562] = t[625] ^ x[35];
  assign t[563] = t[626] ^ x[36];
  assign t[564] = t[627] ^ x[41];
  assign t[565] = t[628] ^ x[42];
  assign t[566] = t[629] ^ x[49];
  assign t[567] = t[630] ^ x[50];
  assign t[568] = t[631] ^ x[55];
  assign t[569] = t[632] ^ x[56];
  assign t[56] = ~(t[89] | t[90]);
  assign t[570] = t[633] ^ x[57];
  assign t[571] = t[634] ^ x[58];
  assign t[572] = t[635] ^ x[63];
  assign t[573] = t[636] ^ x[64];
  assign t[574] = t[637] ^ x[71];
  assign t[575] = t[638] ^ x[72];
  assign t[576] = t[639] ^ x[77];
  assign t[577] = t[640] ^ x[78];
  assign t[578] = t[641] ^ x[79];
  assign t[579] = t[642] ^ x[80];
  assign t[57] = ~(t[91] | t[92]);
  assign t[580] = t[643] ^ x[81];
  assign t[581] = t[644] ^ x[82];
  assign t[582] = t[645] ^ x[83];
  assign t[583] = t[646] ^ x[88];
  assign t[584] = t[647] ^ x[89];
  assign t[585] = t[648] ^ x[92];
  assign t[586] = t[649] ^ x[93];
  assign t[587] = t[650] ^ x[96];
  assign t[588] = t[651] ^ x[97];
  assign t[589] = t[652] ^ x[98];
  assign t[58] = ~(t[413] | t[93]);
  assign t[590] = t[653] ^ x[99];
  assign t[591] = t[654] ^ x[100];
  assign t[592] = t[655] ^ x[103];
  assign t[593] = t[656] ^ x[104];
  assign t[594] = t[657] ^ x[109];
  assign t[595] = t[658] ^ x[110];
  assign t[596] = t[659] ^ x[113];
  assign t[597] = t[660] ^ x[114];
  assign t[598] = t[661] ^ x[115];
  assign t[599] = t[662] ^ x[116];
  assign t[59] = t[30] ? x[44] : x[43];
  assign t[5] = t[9] ^ x[8];
  assign t[600] = t[663] ^ x[117];
  assign t[601] = t[664] ^ x[118];
  assign t[602] = t[665] ^ x[119];
  assign t[603] = t[666] ^ x[120];
  assign t[604] = t[667] ^ x[121];
  assign t[605] = t[668] ^ x[122];
  assign t[606] = t[669] ^ x[123];
  assign t[607] = t[670] ^ x[124];
  assign t[608] = t[671] ^ x[125];
  assign t[609] = t[672] ^ x[141];
  assign t[60] = ~(t[94] & t[95]);
  assign t[610] = t[673] ^ x[157];
  assign t[611] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[612] = (x[0]);
  assign t[613] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[614] = (x[11]);
  assign t[615] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[616] = (x[14]);
  assign t[617] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[618] = (x[17]);
  assign t[619] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = ~(t[96] | t[97]);
  assign t[620] = (x[20]);
  assign t[621] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[622] = (x[24]);
  assign t[623] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[624] = (x[30]);
  assign t[625] = (x[25]);
  assign t[626] = (x[26]);
  assign t[627] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[628] = (x[38]);
  assign t[629] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[62] = ~(t[414] | t[98]);
  assign t[630] = (x[46]);
  assign t[631] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[632] = (x[52]);
  assign t[633] = (x[31]);
  assign t[634] = (x[32]);
  assign t[635] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[636] = (x[60]);
  assign t[637] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[638] = (x[68]);
  assign t[639] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[63] = ~(t[99] | t[100]);
  assign t[640] = (x[74]);
  assign t[641] = (x[23]);
  assign t[642] = (x[39]);
  assign t[643] = (x[40]);
  assign t[644] = (x[47]);
  assign t[645] = (x[48]);
  assign t[646] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[647] = (x[85]);
  assign t[648] = (x[53]);
  assign t[649] = (x[54]);
  assign t[64] = ~(t[101] ^ t[102]);
  assign t[650] = (x[29]);
  assign t[651] = (x[61]);
  assign t[652] = (x[62]);
  assign t[653] = (x[69]);
  assign t[654] = (x[70]);
  assign t[655] = (x[75]);
  assign t[656] = (x[76]);
  assign t[657] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[658] = (x[106]);
  assign t[659] = (x[37]);
  assign t[65] = ~(t[103] | t[104]);
  assign t[660] = (x[45]);
  assign t[661] = (x[86]);
  assign t[662] = (x[87]);
  assign t[663] = (x[51]);
  assign t[664] = (x[59]);
  assign t[665] = (x[67]);
  assign t[666] = (x[73]);
  assign t[667] = (x[107]);
  assign t[668] = (x[108]);
  assign t[669] = (x[84]);
  assign t[66] = ~(t[415] | t[105]);
  assign t[670] = (x[105]);
  assign t[671] = (x[1]);
  assign t[672] = (x[2]);
  assign t[673] = (x[3]);
  assign t[67] = ~(t[106] ^ t[107]);
  assign t[68] = ~(t[416]);
  assign t[69] = ~(t[417]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[110] | t[111]);
  assign t[72] = ~(t[418] | t[112]);
  assign t[73] = t[30] ? x[66] : x[65];
  assign t[74] = ~(t[113] & t[83]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[419] | t[116]);
  assign t[77] = ~(t[117] ^ t[118]);
  assign t[78] = ~(t[119] | t[120]);
  assign t[79] = ~(t[420] | t[121]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[122] | t[123]);
  assign t[81] = ~(t[124] ^ t[125]);
  assign t[82] = ~(t[86] & t[126]);
  assign t[83] = ~(t[127] & t[128]);
  assign t[84] = ~(t[129] | t[130]);
  assign t[85] = ~(t[129] | t[131]);
  assign t[86] = ~(t[132] | t[405]);
  assign t[87] = ~(x[7] | t[406]);
  assign t[88] = x[7] & t[406];
  assign t[89] = ~(t[421]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[411] | t[412]);
  assign t[91] = ~(t[422]);
  assign t[92] = ~(t[423]);
  assign t[93] = ~(t[133] | t[134]);
  assign t[94] = ~(t[135] | t[136]);
  assign t[95] = ~(t[85] | t[137]);
  assign t[96] = ~(t[424]);
  assign t[97] = ~(t[425]);
  assign t[98] = ~(t[138] | t[139]);
  assign t[99] = ~(t[140] | t[141]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[206] & ~t[275] & ~t[354]) | (~t[0] & t[206] & ~t[275] & ~t[354]) | (~t[0] & ~t[206] & t[275] & ~t[354]) | (~t[0] & ~t[206] & ~t[275] & t[354]) | (t[0] & t[206] & t[275] & ~t[354]) | (t[0] & t[206] & ~t[275] & t[354]) | (t[0] & ~t[206] & t[275] & t[354]) | (~t[0] & t[206] & t[275] & t[354]);
endmodule

module R2ind156(x, y);
 input [124:0] x;
 output y;

 wire [364:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[108] | t[98]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[5];
  assign t[156] = t[201] ^ x[13];
  assign t[157] = t[202] ^ x[16];
  assign t[158] = t[203] ^ x[19];
  assign t[159] = t[204] ^ x[22];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[28];
  assign t[161] = t[206] ^ x[36];
  assign t[162] = t[207] ^ x[39];
  assign t[163] = t[208] ^ x[40];
  assign t[164] = t[209] ^ x[46];
  assign t[165] = t[210] ^ x[52];
  assign t[166] = t[211] ^ x[60];
  assign t[167] = t[212] ^ x[63];
  assign t[168] = t[213] ^ x[64];
  assign t[169] = t[214] ^ x[70];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[76];
  assign t[171] = t[216] ^ x[84];
  assign t[172] = t[217] ^ x[87];
  assign t[173] = t[218] ^ x[88];
  assign t[174] = t[219] ^ x[89];
  assign t[175] = t[220] ^ x[90];
  assign t[176] = t[221] ^ x[91];
  assign t[177] = t[222] ^ x[97];
  assign t[178] = t[223] ^ x[98];
  assign t[179] = t[224] ^ x[99];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[100];
  assign t[181] = t[226] ^ x[101];
  assign t[182] = t[227] ^ x[102];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[104];
  assign t[185] = t[230] ^ x[105];
  assign t[186] = t[231] ^ x[106];
  assign t[187] = t[232] ^ x[112];
  assign t[188] = t[233] ^ x[113];
  assign t[189] = t[234] ^ x[114];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[115];
  assign t[191] = t[236] ^ x[116];
  assign t[192] = t[237] ^ x[117];
  assign t[193] = t[238] ^ x[118];
  assign t[194] = t[239] ^ x[119];
  assign t[195] = t[240] ^ x[120];
  assign t[196] = t[241] ^ x[121];
  assign t[197] = t[242] ^ x[122];
  assign t[198] = t[243] ^ x[123];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[245] & t[246]);
  assign t[201] = (~t[247] & t[248]);
  assign t[202] = (~t[249] & t[250]);
  assign t[203] = (~t[251] & t[252]);
  assign t[204] = (~t[253] & t[254]);
  assign t[205] = (~t[255] & t[256]);
  assign t[206] = (~t[257] & t[258]);
  assign t[207] = (~t[255] & t[259]);
  assign t[208] = (~t[255] & t[260]);
  assign t[209] = (~t[261] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[263] & t[264]);
  assign t[211] = (~t[265] & t[266]);
  assign t[212] = (~t[257] & t[267]);
  assign t[213] = (~t[257] & t[268]);
  assign t[214] = (~t[269] & t[270]);
  assign t[215] = (~t[271] & t[272]);
  assign t[216] = (~t[273] & t[274]);
  assign t[217] = (~t[255] & t[275]);
  assign t[218] = (~t[261] & t[276]);
  assign t[219] = (~t[261] & t[277]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[263] & t[278]);
  assign t[221] = (~t[263] & t[279]);
  assign t[222] = (~t[280] & t[281]);
  assign t[223] = (~t[265] & t[282]);
  assign t[224] = (~t[265] & t[283]);
  assign t[225] = (~t[257] & t[284]);
  assign t[226] = (~t[269] & t[285]);
  assign t[227] = (~t[269] & t[286]);
  assign t[228] = (~t[271] & t[287]);
  assign t[229] = (~t[271] & t[288]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[273] & t[289]);
  assign t[231] = (~t[273] & t[290]);
  assign t[232] = (~t[291] & t[292]);
  assign t[233] = (~t[261] & t[293]);
  assign t[234] = (~t[263] & t[294]);
  assign t[235] = (~t[280] & t[295]);
  assign t[236] = (~t[280] & t[296]);
  assign t[237] = (~t[265] & t[297]);
  assign t[238] = (~t[269] & t[298]);
  assign t[239] = (~t[271] & t[299]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[273] & t[300]);
  assign t[241] = (~t[291] & t[301]);
  assign t[242] = (~t[291] & t[302]);
  assign t[243] = (~t[280] & t[303]);
  assign t[244] = (~t[291] & t[304]);
  assign t[245] = t[305] ^ x[4];
  assign t[246] = t[306] ^ x[5];
  assign t[247] = t[307] ^ x[12];
  assign t[248] = t[308] ^ x[13];
  assign t[249] = t[309] ^ x[15];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[310] ^ x[16];
  assign t[251] = t[311] ^ x[18];
  assign t[252] = t[312] ^ x[19];
  assign t[253] = t[313] ^ x[21];
  assign t[254] = t[314] ^ x[22];
  assign t[255] = t[315] ^ x[27];
  assign t[256] = t[316] ^ x[28];
  assign t[257] = t[317] ^ x[35];
  assign t[258] = t[318] ^ x[36];
  assign t[259] = t[319] ^ x[39];
  assign t[25] = ~(t[113]);
  assign t[260] = t[320] ^ x[40];
  assign t[261] = t[321] ^ x[45];
  assign t[262] = t[322] ^ x[46];
  assign t[263] = t[323] ^ x[51];
  assign t[264] = t[324] ^ x[52];
  assign t[265] = t[325] ^ x[59];
  assign t[266] = t[326] ^ x[60];
  assign t[267] = t[327] ^ x[63];
  assign t[268] = t[328] ^ x[64];
  assign t[269] = t[329] ^ x[69];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[70];
  assign t[271] = t[331] ^ x[75];
  assign t[272] = t[332] ^ x[76];
  assign t[273] = t[333] ^ x[83];
  assign t[274] = t[334] ^ x[84];
  assign t[275] = t[335] ^ x[87];
  assign t[276] = t[336] ^ x[88];
  assign t[277] = t[337] ^ x[89];
  assign t[278] = t[338] ^ x[90];
  assign t[279] = t[339] ^ x[91];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[96];
  assign t[281] = t[341] ^ x[97];
  assign t[282] = t[342] ^ x[98];
  assign t[283] = t[343] ^ x[99];
  assign t[284] = t[344] ^ x[100];
  assign t[285] = t[345] ^ x[101];
  assign t[286] = t[346] ^ x[102];
  assign t[287] = t[347] ^ x[103];
  assign t[288] = t[348] ^ x[104];
  assign t[289] = t[349] ^ x[105];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[106];
  assign t[291] = t[351] ^ x[111];
  assign t[292] = t[352] ^ x[112];
  assign t[293] = t[353] ^ x[113];
  assign t[294] = t[354] ^ x[114];
  assign t[295] = t[355] ^ x[115];
  assign t[296] = t[356] ^ x[116];
  assign t[297] = t[357] ^ x[117];
  assign t[298] = t[358] ^ x[118];
  assign t[299] = t[359] ^ x[119];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[120];
  assign t[301] = t[361] ^ x[121];
  assign t[302] = t[362] ^ x[122];
  assign t[303] = t[363] ^ x[123];
  assign t[304] = t[364] ^ x[124];
  assign t[305] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[306] = (x[3]);
  assign t[307] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[308] = (x[11]);
  assign t[309] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = (x[14]);
  assign t[311] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[312] = (x[17]);
  assign t[313] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[314] = (x[20]);
  assign t[315] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[316] = (x[24]);
  assign t[317] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[318] = (x[32]);
  assign t[319] = (x[26]);
  assign t[31] = t[48] | t[115];
  assign t[320] = (x[23]);
  assign t[321] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[322] = (x[42]);
  assign t[323] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[324] = (x[48]);
  assign t[325] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[326] = (x[56]);
  assign t[327] = (x[34]);
  assign t[328] = (x[31]);
  assign t[329] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[32] = t[49] ? x[30] : x[29];
  assign t[330] = (x[66]);
  assign t[331] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[332] = (x[72]);
  assign t[333] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[334] = (x[80]);
  assign t[335] = (x[25]);
  assign t[336] = (x[44]);
  assign t[337] = (x[41]);
  assign t[338] = (x[50]);
  assign t[339] = (x[47]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[92] & ~x[93] & ~x[94] & ~x[95]) | (~x[92] & x[93] & ~x[94] & ~x[95]) | (~x[92] & ~x[93] & x[94] & ~x[95]) | (~x[92] & ~x[93] & ~x[94] & x[95]) | (x[92] & x[93] & x[94] & ~x[95]) | (x[92] & x[93] & ~x[94] & x[95]) | (x[92] & ~x[93] & x[94] & x[95]) | (~x[92] & x[93] & x[94] & x[95]);
  assign t[341] = (x[93]);
  assign t[342] = (x[58]);
  assign t[343] = (x[55]);
  assign t[344] = (x[33]);
  assign t[345] = (x[68]);
  assign t[346] = (x[65]);
  assign t[347] = (x[74]);
  assign t[348] = (x[71]);
  assign t[349] = (x[82]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[79]);
  assign t[351] = (x[107] & ~x[108] & ~x[109] & ~x[110]) | (~x[107] & x[108] & ~x[109] & ~x[110]) | (~x[107] & ~x[108] & x[109] & ~x[110]) | (~x[107] & ~x[108] & ~x[109] & x[110]) | (x[107] & x[108] & x[109] & ~x[110]) | (x[107] & x[108] & ~x[109] & x[110]) | (x[107] & ~x[108] & x[109] & x[110]) | (~x[107] & x[108] & x[109] & x[110]);
  assign t[352] = (x[108]);
  assign t[353] = (x[43]);
  assign t[354] = (x[49]);
  assign t[355] = (x[95]);
  assign t[356] = (x[92]);
  assign t[357] = (x[57]);
  assign t[358] = (x[67]);
  assign t[359] = (x[73]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[81]);
  assign t[361] = (x[110]);
  assign t[362] = (x[107]);
  assign t[363] = (x[94]);
  assign t[364] = (x[109]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[37] = t[58] ^ t[34];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = t[61] | t[116];
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[38] : x[37];
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[44];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[71] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[73]);
  assign t[51] = t[74] | t[119];
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = t[77] | t[120];
  assign t[54] = t[18] ? x[54] : x[53];
  assign t[55] = ~(t[78] & t[79]);
  assign t[56] = ~(t[80] & t[81]);
  assign t[57] = t[82] | t[121];
  assign t[58] = t[18] ? x[62] : x[61];
  assign t[59] = ~(t[122]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[123]);
  assign t[61] = ~(t[83] | t[59]);
  assign t[62] = ~(t[84] & t[85]);
  assign t[63] = t[86] | t[124];
  assign t[64] = ~(t[87] & t[88]);
  assign t[65] = t[89] | t[125];
  assign t[66] = t[90] ? x[78] : x[77];
  assign t[67] = ~(t[91] & t[92]);
  assign t[68] = t[93] | t[126];
  assign t[69] = t[90] ? x[86] : x[85];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[94] & t[95]);
  assign t[71] = ~(t[127]);
  assign t[72] = ~(t[128]);
  assign t[73] = ~(t[129]);
  assign t[74] = ~(t[96] | t[72]);
  assign t[75] = ~(t[130]);
  assign t[76] = ~(t[131]);
  assign t[77] = ~(t[97] | t[75]);
  assign t[78] = ~(t[98] & t[99]);
  assign t[79] = t[100] | t[132];
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[133]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[101] | t[80]);
  assign t[83] = ~(t[135]);
  assign t[84] = ~(t[136]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[102] | t[84]);
  assign t[87] = ~(t[138]);
  assign t[88] = ~(t[139]);
  assign t[89] = ~(t[103] | t[87]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[25]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [124:0] x;
 output y;

 wire [373:0] t;
  assign t[0] = t[1] ? t[2] : t[119];
  assign t[100] = ~(t[153]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[155]);
  assign t[103] = ~(t[115] & t[116]);
  assign t[104] = ~(t[143] & t[142]);
  assign t[105] = ~(t[156]);
  assign t[106] = ~(t[146] & t[145]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[148] & t[147]);
  assign t[109] = ~(t[158]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[117] & t[118]);
  assign t[115] = ~(t[155] & t[154]);
  assign t[116] = ~(t[162]);
  assign t[117] = ~(t[161] & t[160]);
  assign t[118] = ~(t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = t[209] ^ x[5];
  assign t[165] = t[210] ^ x[13];
  assign t[166] = t[211] ^ x[16];
  assign t[167] = t[212] ^ x[19];
  assign t[168] = t[213] ^ x[22];
  assign t[169] = t[214] ^ x[28];
  assign t[16] = ~(t[120] & t[121]);
  assign t[170] = t[215] ^ x[36];
  assign t[171] = t[216] ^ x[39];
  assign t[172] = t[217] ^ x[40];
  assign t[173] = t[218] ^ x[46];
  assign t[174] = t[219] ^ x[52];
  assign t[175] = t[220] ^ x[60];
  assign t[176] = t[221] ^ x[63];
  assign t[177] = t[222] ^ x[64];
  assign t[178] = t[223] ^ x[70];
  assign t[179] = t[224] ^ x[76];
  assign t[17] = ~(t[122] & t[123]);
  assign t[180] = t[225] ^ x[84];
  assign t[181] = t[226] ^ x[87];
  assign t[182] = t[227] ^ x[88];
  assign t[183] = t[228] ^ x[89];
  assign t[184] = t[229] ^ x[90];
  assign t[185] = t[230] ^ x[91];
  assign t[186] = t[231] ^ x[97];
  assign t[187] = t[232] ^ x[98];
  assign t[188] = t[233] ^ x[99];
  assign t[189] = t[234] ^ x[100];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[101];
  assign t[191] = t[236] ^ x[102];
  assign t[192] = t[237] ^ x[103];
  assign t[193] = t[238] ^ x[104];
  assign t[194] = t[239] ^ x[105];
  assign t[195] = t[240] ^ x[106];
  assign t[196] = t[241] ^ x[112];
  assign t[197] = t[242] ^ x[113];
  assign t[198] = t[243] ^ x[114];
  assign t[199] = t[244] ^ x[115];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[116];
  assign t[201] = t[246] ^ x[117];
  assign t[202] = t[247] ^ x[118];
  assign t[203] = t[248] ^ x[119];
  assign t[204] = t[249] ^ x[120];
  assign t[205] = t[250] ^ x[121];
  assign t[206] = t[251] ^ x[122];
  assign t[207] = t[252] ^ x[123];
  assign t[208] = t[253] ^ x[124];
  assign t[209] = (~t[254] & t[255]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[256] & t[257]);
  assign t[211] = (~t[258] & t[259]);
  assign t[212] = (~t[260] & t[261]);
  assign t[213] = (~t[262] & t[263]);
  assign t[214] = (~t[264] & t[265]);
  assign t[215] = (~t[266] & t[267]);
  assign t[216] = (~t[264] & t[268]);
  assign t[217] = (~t[264] & t[269]);
  assign t[218] = (~t[270] & t[271]);
  assign t[219] = (~t[272] & t[273]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[274] & t[275]);
  assign t[221] = (~t[266] & t[276]);
  assign t[222] = (~t[266] & t[277]);
  assign t[223] = (~t[278] & t[279]);
  assign t[224] = (~t[280] & t[281]);
  assign t[225] = (~t[282] & t[283]);
  assign t[226] = (~t[264] & t[284]);
  assign t[227] = (~t[270] & t[285]);
  assign t[228] = (~t[270] & t[286]);
  assign t[229] = (~t[272] & t[287]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[272] & t[288]);
  assign t[231] = (~t[289] & t[290]);
  assign t[232] = (~t[274] & t[291]);
  assign t[233] = (~t[274] & t[292]);
  assign t[234] = (~t[266] & t[293]);
  assign t[235] = (~t[278] & t[294]);
  assign t[236] = (~t[278] & t[295]);
  assign t[237] = (~t[280] & t[296]);
  assign t[238] = (~t[280] & t[297]);
  assign t[239] = (~t[282] & t[298]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[282] & t[299]);
  assign t[241] = (~t[300] & t[301]);
  assign t[242] = (~t[270] & t[302]);
  assign t[243] = (~t[272] & t[303]);
  assign t[244] = (~t[289] & t[304]);
  assign t[245] = (~t[289] & t[305]);
  assign t[246] = (~t[274] & t[306]);
  assign t[247] = (~t[278] & t[307]);
  assign t[248] = (~t[280] & t[308]);
  assign t[249] = (~t[282] & t[309]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = (~t[300] & t[310]);
  assign t[251] = (~t[300] & t[311]);
  assign t[252] = (~t[289] & t[312]);
  assign t[253] = (~t[300] & t[313]);
  assign t[254] = t[314] ^ x[4];
  assign t[255] = t[315] ^ x[5];
  assign t[256] = t[316] ^ x[12];
  assign t[257] = t[317] ^ x[13];
  assign t[258] = t[318] ^ x[15];
  assign t[259] = t[319] ^ x[16];
  assign t[25] = ~(t[122]);
  assign t[260] = t[320] ^ x[18];
  assign t[261] = t[321] ^ x[19];
  assign t[262] = t[322] ^ x[21];
  assign t[263] = t[323] ^ x[22];
  assign t[264] = t[324] ^ x[27];
  assign t[265] = t[325] ^ x[28];
  assign t[266] = t[326] ^ x[35];
  assign t[267] = t[327] ^ x[36];
  assign t[268] = t[328] ^ x[39];
  assign t[269] = t[329] ^ x[40];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[45];
  assign t[271] = t[331] ^ x[46];
  assign t[272] = t[332] ^ x[51];
  assign t[273] = t[333] ^ x[52];
  assign t[274] = t[334] ^ x[59];
  assign t[275] = t[335] ^ x[60];
  assign t[276] = t[336] ^ x[63];
  assign t[277] = t[337] ^ x[64];
  assign t[278] = t[338] ^ x[69];
  assign t[279] = t[339] ^ x[70];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[75];
  assign t[281] = t[341] ^ x[76];
  assign t[282] = t[342] ^ x[83];
  assign t[283] = t[343] ^ x[84];
  assign t[284] = t[344] ^ x[87];
  assign t[285] = t[345] ^ x[88];
  assign t[286] = t[346] ^ x[89];
  assign t[287] = t[347] ^ x[90];
  assign t[288] = t[348] ^ x[91];
  assign t[289] = t[349] ^ x[96];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[97];
  assign t[291] = t[351] ^ x[98];
  assign t[292] = t[352] ^ x[99];
  assign t[293] = t[353] ^ x[100];
  assign t[294] = t[354] ^ x[101];
  assign t[295] = t[355] ^ x[102];
  assign t[296] = t[356] ^ x[103];
  assign t[297] = t[357] ^ x[104];
  assign t[298] = t[358] ^ x[105];
  assign t[299] = t[359] ^ x[106];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[111];
  assign t[301] = t[361] ^ x[112];
  assign t[302] = t[362] ^ x[113];
  assign t[303] = t[363] ^ x[114];
  assign t[304] = t[364] ^ x[115];
  assign t[305] = t[365] ^ x[116];
  assign t[306] = t[366] ^ x[117];
  assign t[307] = t[367] ^ x[118];
  assign t[308] = t[368] ^ x[119];
  assign t[309] = t[369] ^ x[120];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[370] ^ x[121];
  assign t[311] = t[371] ^ x[122];
  assign t[312] = t[372] ^ x[123];
  assign t[313] = t[373] ^ x[124];
  assign t[314] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[315] = (x[2]);
  assign t[316] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[317] = (x[11]);
  assign t[318] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[319] = (x[14]);
  assign t[31] = ~(t[48] & t[124]);
  assign t[320] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[321] = (x[17]);
  assign t[322] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[323] = (x[20]);
  assign t[324] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[325] = (x[24]);
  assign t[326] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[327] = (x[32]);
  assign t[328] = (x[26]);
  assign t[329] = (x[23]);
  assign t[32] = t[49] ? x[30] : x[29];
  assign t[330] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[331] = (x[42]);
  assign t[332] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[333] = (x[48]);
  assign t[334] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[335] = (x[56]);
  assign t[336] = (x[34]);
  assign t[337] = (x[31]);
  assign t[338] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[339] = (x[66]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[341] = (x[72]);
  assign t[342] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[343] = (x[80]);
  assign t[344] = (x[25]);
  assign t[345] = (x[44]);
  assign t[346] = (x[41]);
  assign t[347] = (x[50]);
  assign t[348] = (x[47]);
  assign t[349] = (x[92] & ~x[93] & ~x[94] & ~x[95]) | (~x[92] & x[93] & ~x[94] & ~x[95]) | (~x[92] & ~x[93] & x[94] & ~x[95]) | (~x[92] & ~x[93] & ~x[94] & x[95]) | (x[92] & x[93] & x[94] & ~x[95]) | (x[92] & x[93] & ~x[94] & x[95]) | (x[92] & ~x[93] & x[94] & x[95]) | (~x[92] & x[93] & x[94] & x[95]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[93]);
  assign t[351] = (x[58]);
  assign t[352] = (x[55]);
  assign t[353] = (x[33]);
  assign t[354] = (x[68]);
  assign t[355] = (x[65]);
  assign t[356] = (x[74]);
  assign t[357] = (x[71]);
  assign t[358] = (x[82]);
  assign t[359] = (x[79]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[107] & ~x[108] & ~x[109] & ~x[110]) | (~x[107] & x[108] & ~x[109] & ~x[110]) | (~x[107] & ~x[108] & x[109] & ~x[110]) | (~x[107] & ~x[108] & ~x[109] & x[110]) | (x[107] & x[108] & x[109] & ~x[110]) | (x[107] & x[108] & ~x[109] & x[110]) | (x[107] & ~x[108] & x[109] & x[110]) | (~x[107] & x[108] & x[109] & x[110]);
  assign t[361] = (x[108]);
  assign t[362] = (x[43]);
  assign t[363] = (x[49]);
  assign t[364] = (x[95]);
  assign t[365] = (x[92]);
  assign t[366] = (x[57]);
  assign t[367] = (x[67]);
  assign t[368] = (x[73]);
  assign t[369] = (x[81]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[110]);
  assign t[371] = (x[107]);
  assign t[372] = (x[94]);
  assign t[373] = (x[109]);
  assign t[37] = t[58] ^ t[34];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = ~(t[61] & t[125]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[38] : x[37];
  assign t[41] = ~(t[62] & t[63]);
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[44];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[70];
  assign t[46] = ~(t[126]);
  assign t[47] = ~(t[127]);
  assign t[48] = ~(t[71] & t[72]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = ~(t[75] & t[128]);
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = ~(t[78] & t[129]);
  assign t[54] = t[18] ? x[54] : x[53];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = ~(t[83] & t[130]);
  assign t[58] = t[122] ? x[62] : x[61];
  assign t[59] = ~(t[131]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[132]);
  assign t[61] = ~(t[84] & t[85]);
  assign t[62] = ~(t[86] & t[87]);
  assign t[63] = ~(t[88] & t[133]);
  assign t[64] = ~(t[89] & t[90]);
  assign t[65] = ~(t[91] & t[134]);
  assign t[66] = t[49] ? x[78] : x[77];
  assign t[67] = ~(t[92] & t[93]);
  assign t[68] = ~(t[94] & t[135]);
  assign t[69] = t[49] ? x[86] : x[85];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[95] & t[96]);
  assign t[71] = ~(t[127] & t[126]);
  assign t[72] = ~(t[136]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[97] & t[98]);
  assign t[76] = ~(t[139]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[99] & t[100]);
  assign t[79] = ~(t[101] & t[102]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[103] & t[141]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[104] & t[105]);
  assign t[84] = ~(t[132] & t[131]);
  assign t[85] = ~(t[144]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[106] & t[107]);
  assign t[89] = ~(t[147]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[108] & t[109]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[150]);
  assign t[94] = ~(t[110] & t[111]);
  assign t[95] = ~(t[112] & t[113]);
  assign t[96] = ~(t[114] & t[151]);
  assign t[97] = ~(t[138] & t[137]);
  assign t[98] = ~(t[152]);
  assign t[99] = ~(t[140] & t[139]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [114:0] x;
 output y;

 wire [303:0] t;
  assign t[0] = t[1] ? t[2] : t[99];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = t[169] ^ x[5];
  assign t[135] = t[170] ^ x[13];
  assign t[136] = t[171] ^ x[16];
  assign t[137] = t[172] ^ x[19];
  assign t[138] = t[173] ^ x[22];
  assign t[139] = t[174] ^ x[28];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[29];
  assign t[141] = t[176] ^ x[37];
  assign t[142] = t[177] ^ x[38];
  assign t[143] = t[178] ^ x[41];
  assign t[144] = t[179] ^ x[47];
  assign t[145] = t[180] ^ x[48];
  assign t[146] = t[181] ^ x[54];
  assign t[147] = t[182] ^ x[55];
  assign t[148] = t[183] ^ x[63];
  assign t[149] = t[184] ^ x[64];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[67];
  assign t[151] = t[186] ^ x[73];
  assign t[152] = t[187] ^ x[74];
  assign t[153] = t[188] ^ x[80];
  assign t[154] = t[189] ^ x[81];
  assign t[155] = t[190] ^ x[89];
  assign t[156] = t[191] ^ x[90];
  assign t[157] = t[192] ^ x[93];
  assign t[158] = t[193] ^ x[94];
  assign t[159] = t[194] ^ x[95];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[101];
  assign t[161] = t[196] ^ x[102];
  assign t[162] = t[197] ^ x[103];
  assign t[163] = t[198] ^ x[104];
  assign t[164] = t[199] ^ x[110];
  assign t[165] = t[200] ^ x[111];
  assign t[166] = t[201] ^ x[112];
  assign t[167] = t[202] ^ x[113];
  assign t[168] = t[203] ^ x[114];
  assign t[169] = (~t[204] & t[205]);
  assign t[16] = ~(t[100] & t[101]);
  assign t[170] = (~t[206] & t[207]);
  assign t[171] = (~t[208] & t[209]);
  assign t[172] = (~t[210] & t[211]);
  assign t[173] = (~t[212] & t[213]);
  assign t[174] = (~t[214] & t[215]);
  assign t[175] = (~t[214] & t[216]);
  assign t[176] = (~t[217] & t[218]);
  assign t[177] = (~t[217] & t[219]);
  assign t[178] = (~t[214] & t[220]);
  assign t[179] = (~t[221] & t[222]);
  assign t[17] = ~(t[102] & t[103]);
  assign t[180] = (~t[221] & t[223]);
  assign t[181] = (~t[224] & t[225]);
  assign t[182] = (~t[224] & t[226]);
  assign t[183] = (~t[227] & t[228]);
  assign t[184] = (~t[227] & t[229]);
  assign t[185] = (~t[217] & t[230]);
  assign t[186] = (~t[231] & t[232]);
  assign t[187] = (~t[231] & t[233]);
  assign t[188] = (~t[234] & t[235]);
  assign t[189] = (~t[234] & t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (~t[237] & t[238]);
  assign t[191] = (~t[237] & t[239]);
  assign t[192] = (~t[221] & t[240]);
  assign t[193] = (~t[224] & t[241]);
  assign t[194] = (~t[227] & t[242]);
  assign t[195] = (~t[243] & t[244]);
  assign t[196] = (~t[243] & t[245]);
  assign t[197] = (~t[231] & t[246]);
  assign t[198] = (~t[234] & t[247]);
  assign t[199] = (~t[248] & t[249]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[248] & t[250]);
  assign t[201] = (~t[237] & t[251]);
  assign t[202] = (~t[243] & t[252]);
  assign t[203] = (~t[248] & t[253]);
  assign t[204] = t[254] ^ x[4];
  assign t[205] = t[255] ^ x[5];
  assign t[206] = t[256] ^ x[12];
  assign t[207] = t[257] ^ x[13];
  assign t[208] = t[258] ^ x[15];
  assign t[209] = t[259] ^ x[16];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[260] ^ x[18];
  assign t[211] = t[261] ^ x[19];
  assign t[212] = t[262] ^ x[21];
  assign t[213] = t[263] ^ x[22];
  assign t[214] = t[264] ^ x[27];
  assign t[215] = t[265] ^ x[28];
  assign t[216] = t[266] ^ x[29];
  assign t[217] = t[267] ^ x[36];
  assign t[218] = t[268] ^ x[37];
  assign t[219] = t[269] ^ x[38];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[270] ^ x[41];
  assign t[221] = t[271] ^ x[46];
  assign t[222] = t[272] ^ x[47];
  assign t[223] = t[273] ^ x[48];
  assign t[224] = t[274] ^ x[53];
  assign t[225] = t[275] ^ x[54];
  assign t[226] = t[276] ^ x[55];
  assign t[227] = t[277] ^ x[62];
  assign t[228] = t[278] ^ x[63];
  assign t[229] = t[279] ^ x[64];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[280] ^ x[67];
  assign t[231] = t[281] ^ x[72];
  assign t[232] = t[282] ^ x[73];
  assign t[233] = t[283] ^ x[74];
  assign t[234] = t[284] ^ x[79];
  assign t[235] = t[285] ^ x[80];
  assign t[236] = t[286] ^ x[81];
  assign t[237] = t[287] ^ x[88];
  assign t[238] = t[288] ^ x[89];
  assign t[239] = t[289] ^ x[90];
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = t[290] ^ x[93];
  assign t[241] = t[291] ^ x[94];
  assign t[242] = t[292] ^ x[95];
  assign t[243] = t[293] ^ x[100];
  assign t[244] = t[294] ^ x[101];
  assign t[245] = t[295] ^ x[102];
  assign t[246] = t[296] ^ x[103];
  assign t[247] = t[297] ^ x[104];
  assign t[248] = t[298] ^ x[109];
  assign t[249] = t[299] ^ x[110];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[300] ^ x[111];
  assign t[251] = t[301] ^ x[112];
  assign t[252] = t[302] ^ x[113];
  assign t[253] = t[303] ^ x[114];
  assign t[254] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[255] = (x[1]);
  assign t[256] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[257] = (x[11]);
  assign t[258] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[259] = (x[14]);
  assign t[25] = ~(t[102]);
  assign t[260] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[261] = (x[17]);
  assign t[262] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[263] = (x[20]);
  assign t[264] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[265] = (x[25]);
  assign t[266] = (x[23]);
  assign t[267] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[268] = (x[34]);
  assign t[269] = (x[32]);
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = (x[26]);
  assign t[271] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[272] = (x[44]);
  assign t[273] = (x[42]);
  assign t[274] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[275] = (x[51]);
  assign t[276] = (x[49]);
  assign t[277] = (x[58] & ~x[59] & ~x[60] & ~x[61]) | (~x[58] & x[59] & ~x[60] & ~x[61]) | (~x[58] & ~x[59] & x[60] & ~x[61]) | (~x[58] & ~x[59] & ~x[60] & x[61]) | (x[58] & x[59] & x[60] & ~x[61]) | (x[58] & x[59] & ~x[60] & x[61]) | (x[58] & ~x[59] & x[60] & x[61]) | (~x[58] & x[59] & x[60] & x[61]);
  assign t[278] = (x[60]);
  assign t[279] = (x[58]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[35]);
  assign t[281] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[282] = (x[70]);
  assign t[283] = (x[68]);
  assign t[284] = (x[75] & ~x[76] & ~x[77] & ~x[78]) | (~x[75] & x[76] & ~x[77] & ~x[78]) | (~x[75] & ~x[76] & x[77] & ~x[78]) | (~x[75] & ~x[76] & ~x[77] & x[78]) | (x[75] & x[76] & x[77] & ~x[78]) | (x[75] & x[76] & ~x[77] & x[78]) | (x[75] & ~x[76] & x[77] & x[78]) | (~x[75] & x[76] & x[77] & x[78]);
  assign t[285] = (x[77]);
  assign t[286] = (x[75]);
  assign t[287] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[288] = (x[86]);
  assign t[289] = (x[84]);
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = (x[45]);
  assign t[291] = (x[52]);
  assign t[292] = (x[61]);
  assign t[293] = (x[96] & ~x[97] & ~x[98] & ~x[99]) | (~x[96] & x[97] & ~x[98] & ~x[99]) | (~x[96] & ~x[97] & x[98] & ~x[99]) | (~x[96] & ~x[97] & ~x[98] & x[99]) | (x[96] & x[97] & x[98] & ~x[99]) | (x[96] & x[97] & ~x[98] & x[99]) | (x[96] & ~x[97] & x[98] & x[99]) | (~x[96] & x[97] & x[98] & x[99]);
  assign t[294] = (x[98]);
  assign t[295] = (x[96]);
  assign t[296] = (x[71]);
  assign t[297] = (x[78]);
  assign t[298] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[299] = (x[107]);
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[105]);
  assign t[301] = (x[87]);
  assign t[302] = (x[99]);
  assign t[303] = (x[108]);
  assign t[30] = ~(t[104] & t[46]);
  assign t[31] = ~(t[105] & t[47]);
  assign t[32] = t[18] ? x[31] : x[30];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[36];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = t[55] ^ t[56];
  assign t[38] = ~(t[106] & t[57]);
  assign t[39] = ~(t[107] & t[58]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[40] : x[39];
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = ~(t[61] & t[62]);
  assign t[43] = t[63] ^ t[64];
  assign t[44] = ~(t[65] & t[66]);
  assign t[45] = t[67] ^ t[42];
  assign t[46] = ~(t[108]);
  assign t[47] = ~(t[108] & t[68]);
  assign t[48] = ~(t[109] & t[69]);
  assign t[49] = ~(t[110] & t[70]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[71]);
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = t[73] ? x[57] : x[56];
  assign t[53] = ~(t[113] & t[74]);
  assign t[54] = ~(t[114] & t[75]);
  assign t[55] = t[18] ? x[66] : x[65];
  assign t[56] = ~(t[76] & t[77]);
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[115] & t[78]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[117] & t[80]);
  assign t[61] = ~(t[118] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = t[73] ? x[83] : x[82];
  assign t[64] = ~(t[83] & t[84]);
  assign t[65] = ~(t[120] & t[85]);
  assign t[66] = ~(t[121] & t[86]);
  assign t[67] = t[73] ? x[92] : x[91];
  assign t[68] = ~(t[104]);
  assign t[69] = ~(t[122]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[122] & t[87]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[25]);
  assign t[74] = ~(t[124]);
  assign t[75] = ~(t[124] & t[89]);
  assign t[76] = ~(t[125] & t[90]);
  assign t[77] = ~(t[126] & t[91]);
  assign t[78] = ~(t[106]);
  assign t[79] = ~(t[127]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127] & t[92]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[128] & t[93]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130] & t[95]);
  assign t[85] = ~(t[131]);
  assign t[86] = ~(t[131] & t[96]);
  assign t[87] = ~(t[109]);
  assign t[88] = ~(t[111]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[132]);
  assign t[91] = ~(t[132] & t[97]);
  assign t[92] = ~(t[116]);
  assign t[93] = ~(t[118]);
  assign t[94] = ~(t[133]);
  assign t[95] = ~(t[133] & t[98]);
  assign t[96] = ~(t[120]);
  assign t[97] = ~(t[125]);
  assign t[98] = ~(t[129]);
  assign t[99] = (t[134]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [124:0] x;
 output y;

 wire [460:0] t;
  assign t[0] = t[1] ? t[2] : t[206];
  assign t[100] = ~(t[228] | t[142]);
  assign t[101] = t[30] ? x[91] : x[90];
  assign t[102] = ~(t[143] & t[144]);
  assign t[103] = ~(t[229]);
  assign t[104] = ~(t[230]);
  assign t[105] = ~(t[145] | t[146]);
  assign t[106] = t[30] ? x[95] : x[94];
  assign t[107] = ~(t[147] & t[148]);
  assign t[108] = ~(t[231]);
  assign t[109] = ~(t[218] | t[219]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[232]);
  assign t[111] = ~(t[233]);
  assign t[112] = ~(t[149] | t[150]);
  assign t[113] = ~(t[151] | t[152]);
  assign t[114] = ~(t[234]);
  assign t[115] = ~(t[235]);
  assign t[116] = ~(t[153] | t[154]);
  assign t[117] = t[155] ? x[102] : x[101];
  assign t[118] = t[156] | t[84];
  assign t[119] = ~(t[236]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[237]);
  assign t[121] = ~(t[157] | t[158]);
  assign t[122] = ~(t[159] | t[160]);
  assign t[123] = ~(t[238] | t[161]);
  assign t[124] = t[155] ? x[112] : x[111];
  assign t[125] = ~(t[162] & t[163]);
  assign t[126] = ~(t[164] & t[165]);
  assign t[127] = ~(t[208] | t[166]);
  assign t[128] = t[129] & t[207];
  assign t[129] = ~(t[132]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[207] ? t[164] : t[167];
  assign t[131] = t[207] ? t[169] : t[168];
  assign t[132] = ~(t[209]);
  assign t[133] = ~(t[239]);
  assign t[134] = ~(t[224] | t[225]);
  assign t[135] = ~(t[132] | t[170]);
  assign t[136] = ~(t[129] | t[171]);
  assign t[137] = ~(t[172] & t[173]);
  assign t[138] = ~(t[240]);
  assign t[139] = ~(t[226] | t[227]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[241]);
  assign t[141] = ~(t[242]);
  assign t[142] = ~(t[174] | t[175]);
  assign t[143] = ~(t[151] | t[176]);
  assign t[144] = ~(t[118] | t[177]);
  assign t[145] = ~(t[243]);
  assign t[146] = ~(t[229] | t[230]);
  assign t[147] = ~(t[178] | t[85]);
  assign t[148] = ~(t[135] | t[156]);
  assign t[149] = ~(t[244]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[232] | t[233]);
  assign t[151] = ~(t[129] | t[179]);
  assign t[152] = ~(t[94] & t[180]);
  assign t[153] = ~(t[245]);
  assign t[154] = ~(t[234] | t[235]);
  assign t[155] = ~(t[49]);
  assign t[156] = ~(t[181] & t[83]);
  assign t[157] = ~(t[246]);
  assign t[158] = ~(t[236] | t[237]);
  assign t[159] = ~(t[247]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[248]);
  assign t[161] = ~(t[182] | t[183]);
  assign t[162] = ~(t[151]);
  assign t[163] = ~(t[184] | t[84]);
  assign t[164] = ~(t[210] & t[185]);
  assign t[165] = ~(x[7] & t[127]);
  assign t[166] = ~(t[210]);
  assign t[167] = ~(x[7] & t[186]);
  assign t[168] = ~(t[88] & t[166]);
  assign t[169] = ~(t[87] & t[210]);
  assign t[16] = ~(t[207] & t[208]);
  assign t[170] = t[207] ? t[187] : t[168];
  assign t[171] = t[207] ? t[188] : t[165];
  assign t[172] = ~(t[151] | t[189]);
  assign t[173] = t[132] | t[190];
  assign t[174] = ~(t[249]);
  assign t[175] = ~(t[241] | t[242]);
  assign t[176] = ~(t[129] | t[191]);
  assign t[177] = ~(t[192] & t[173]);
  assign t[178] = ~(t[129] | t[193]);
  assign t[179] = t[207] ? t[194] : t[187];
  assign t[17] = ~(t[209] & t[210]);
  assign t[180] = ~(t[132] & t[195]);
  assign t[181] = ~(t[196] | t[197]);
  assign t[182] = ~(t[250]);
  assign t[183] = ~(t[247] | t[248]);
  assign t[184] = ~(t[198]);
  assign t[185] = ~(x[7] | t[199]);
  assign t[186] = ~(t[208] | t[210]);
  assign t[187] = ~(t[87] & t[166]);
  assign t[188] = ~(t[185] & t[166]);
  assign t[189] = ~(t[129] | t[200]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = t[207] ? t[167] : t[188];
  assign t[191] = t[207] ? t[167] : t[164];
  assign t[192] = ~(t[201] | t[202]);
  assign t[193] = t[207] ? t[187] : t[194];
  assign t[194] = ~(t[88] & t[210]);
  assign t[195] = ~(t[167] & t[164]);
  assign t[196] = ~(t[132] | t[203]);
  assign t[197] = ~(t[132] | t[204]);
  assign t[198] = ~(t[202] | t[189]);
  assign t[199] = ~(t[208]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[207] ? t[168] : t[169];
  assign t[201] = ~(t[82]);
  assign t[202] = ~(t[129] | t[205]);
  assign t[203] = t[207] ? t[168] : t[187];
  assign t[204] = t[207] ? t[188] : t[167];
  assign t[205] = t[207] ? t[165] : t[188];
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = t[296] ^ x[5];
  assign t[252] = t[297] ^ x[13];
  assign t[253] = t[298] ^ x[16];
  assign t[254] = t[299] ^ x[19];
  assign t[255] = t[300] ^ x[22];
  assign t[256] = t[301] ^ x[28];
  assign t[257] = t[302] ^ x[34];
  assign t[258] = t[303] ^ x[35];
  assign t[259] = t[304] ^ x[36];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[42];
  assign t[261] = t[306] ^ x[50];
  assign t[262] = t[307] ^ x[56];
  assign t[263] = t[308] ^ x[57];
  assign t[264] = t[309] ^ x[58];
  assign t[265] = t[310] ^ x[64];
  assign t[266] = t[311] ^ x[72];
  assign t[267] = t[312] ^ x[78];
  assign t[268] = t[313] ^ x[79];
  assign t[269] = t[314] ^ x[80];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[81];
  assign t[271] = t[316] ^ x[82];
  assign t[272] = t[317] ^ x[83];
  assign t[273] = t[318] ^ x[89];
  assign t[274] = t[319] ^ x[92];
  assign t[275] = t[320] ^ x[93];
  assign t[276] = t[321] ^ x[96];
  assign t[277] = t[322] ^ x[97];
  assign t[278] = t[323] ^ x[98];
  assign t[279] = t[324] ^ x[99];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[100];
  assign t[281] = t[326] ^ x[103];
  assign t[282] = t[327] ^ x[104];
  assign t[283] = t[328] ^ x[110];
  assign t[284] = t[329] ^ x[113];
  assign t[285] = t[330] ^ x[114];
  assign t[286] = t[331] ^ x[115];
  assign t[287] = t[332] ^ x[116];
  assign t[288] = t[333] ^ x[117];
  assign t[289] = t[334] ^ x[118];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[119];
  assign t[291] = t[336] ^ x[120];
  assign t[292] = t[337] ^ x[121];
  assign t[293] = t[338] ^ x[122];
  assign t[294] = t[339] ^ x[123];
  assign t[295] = t[340] ^ x[124];
  assign t[296] = (~t[341] & t[342]);
  assign t[297] = (~t[343] & t[344]);
  assign t[298] = (~t[345] & t[346]);
  assign t[299] = (~t[347] & t[348]);
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[349] & t[350]);
  assign t[301] = (~t[351] & t[352]);
  assign t[302] = (~t[353] & t[354]);
  assign t[303] = (~t[351] & t[355]);
  assign t[304] = (~t[351] & t[356]);
  assign t[305] = (~t[357] & t[358]);
  assign t[306] = (~t[359] & t[360]);
  assign t[307] = (~t[361] & t[362]);
  assign t[308] = (~t[353] & t[363]);
  assign t[309] = (~t[353] & t[364]);
  assign t[30] = ~(t[49]);
  assign t[310] = (~t[365] & t[366]);
  assign t[311] = (~t[367] & t[368]);
  assign t[312] = (~t[369] & t[370]);
  assign t[313] = (~t[351] & t[371]);
  assign t[314] = (~t[357] & t[372]);
  assign t[315] = (~t[357] & t[373]);
  assign t[316] = (~t[359] & t[374]);
  assign t[317] = (~t[359] & t[375]);
  assign t[318] = (~t[376] & t[377]);
  assign t[319] = (~t[361] & t[378]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (~t[361] & t[379]);
  assign t[321] = (~t[353] & t[380]);
  assign t[322] = (~t[365] & t[381]);
  assign t[323] = (~t[365] & t[382]);
  assign t[324] = (~t[367] & t[383]);
  assign t[325] = (~t[367] & t[384]);
  assign t[326] = (~t[369] & t[385]);
  assign t[327] = (~t[369] & t[386]);
  assign t[328] = (~t[387] & t[388]);
  assign t[329] = (~t[357] & t[389]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[330] = (~t[359] & t[390]);
  assign t[331] = (~t[376] & t[391]);
  assign t[332] = (~t[376] & t[392]);
  assign t[333] = (~t[361] & t[393]);
  assign t[334] = (~t[365] & t[394]);
  assign t[335] = (~t[367] & t[395]);
  assign t[336] = (~t[369] & t[396]);
  assign t[337] = (~t[387] & t[397]);
  assign t[338] = (~t[387] & t[398]);
  assign t[339] = (~t[376] & t[399]);
  assign t[33] = ~(t[54] | t[55]);
  assign t[340] = (~t[387] & t[400]);
  assign t[341] = t[401] ^ x[4];
  assign t[342] = t[402] ^ x[5];
  assign t[343] = t[403] ^ x[12];
  assign t[344] = t[404] ^ x[13];
  assign t[345] = t[405] ^ x[15];
  assign t[346] = t[406] ^ x[16];
  assign t[347] = t[407] ^ x[18];
  assign t[348] = t[408] ^ x[19];
  assign t[349] = t[409] ^ x[21];
  assign t[34] = ~(t[211] | t[56]);
  assign t[350] = t[410] ^ x[22];
  assign t[351] = t[411] ^ x[27];
  assign t[352] = t[412] ^ x[28];
  assign t[353] = t[413] ^ x[33];
  assign t[354] = t[414] ^ x[34];
  assign t[355] = t[415] ^ x[35];
  assign t[356] = t[416] ^ x[36];
  assign t[357] = t[417] ^ x[41];
  assign t[358] = t[418] ^ x[42];
  assign t[359] = t[419] ^ x[49];
  assign t[35] = ~(t[57] | t[58]);
  assign t[360] = t[420] ^ x[50];
  assign t[361] = t[421] ^ x[55];
  assign t[362] = t[422] ^ x[56];
  assign t[363] = t[423] ^ x[57];
  assign t[364] = t[424] ^ x[58];
  assign t[365] = t[425] ^ x[63];
  assign t[366] = t[426] ^ x[64];
  assign t[367] = t[427] ^ x[71];
  assign t[368] = t[428] ^ x[72];
  assign t[369] = t[429] ^ x[77];
  assign t[36] = ~(t[59] ^ t[60]);
  assign t[370] = t[430] ^ x[78];
  assign t[371] = t[431] ^ x[79];
  assign t[372] = t[432] ^ x[80];
  assign t[373] = t[433] ^ x[81];
  assign t[374] = t[434] ^ x[82];
  assign t[375] = t[435] ^ x[83];
  assign t[376] = t[436] ^ x[88];
  assign t[377] = t[437] ^ x[89];
  assign t[378] = t[438] ^ x[92];
  assign t[379] = t[439] ^ x[93];
  assign t[37] = ~(t[61] | t[62]);
  assign t[380] = t[440] ^ x[96];
  assign t[381] = t[441] ^ x[97];
  assign t[382] = t[442] ^ x[98];
  assign t[383] = t[443] ^ x[99];
  assign t[384] = t[444] ^ x[100];
  assign t[385] = t[445] ^ x[103];
  assign t[386] = t[446] ^ x[104];
  assign t[387] = t[447] ^ x[109];
  assign t[388] = t[448] ^ x[110];
  assign t[389] = t[449] ^ x[113];
  assign t[38] = ~(t[63] ^ t[64]);
  assign t[390] = t[450] ^ x[114];
  assign t[391] = t[451] ^ x[115];
  assign t[392] = t[452] ^ x[116];
  assign t[393] = t[453] ^ x[117];
  assign t[394] = t[454] ^ x[118];
  assign t[395] = t[455] ^ x[119];
  assign t[396] = t[456] ^ x[120];
  assign t[397] = t[457] ^ x[121];
  assign t[398] = t[458] ^ x[122];
  assign t[399] = t[459] ^ x[123];
  assign t[39] = ~(t[65] | t[66]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[460] ^ x[124];
  assign t[401] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[402] = (x[0]);
  assign t[403] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[404] = (x[11]);
  assign t[405] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[406] = (x[14]);
  assign t[407] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[408] = (x[17]);
  assign t[409] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[40] = ~(t[37] ^ t[67]);
  assign t[410] = (x[20]);
  assign t[411] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[412] = (x[24]);
  assign t[413] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[414] = (x[30]);
  assign t[415] = (x[25]);
  assign t[416] = (x[26]);
  assign t[417] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[418] = (x[38]);
  assign t[419] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[41] = ~(t[68] | t[69]);
  assign t[420] = (x[46]);
  assign t[421] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[422] = (x[52]);
  assign t[423] = (x[31]);
  assign t[424] = (x[32]);
  assign t[425] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[426] = (x[60]);
  assign t[427] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[428] = (x[68]);
  assign t[429] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[42] = ~(t[212] | t[70]);
  assign t[430] = (x[74]);
  assign t[431] = (x[23]);
  assign t[432] = (x[39]);
  assign t[433] = (x[40]);
  assign t[434] = (x[47]);
  assign t[435] = (x[48]);
  assign t[436] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[437] = (x[85]);
  assign t[438] = (x[53]);
  assign t[439] = (x[54]);
  assign t[43] = ~(t[71] | t[72]);
  assign t[440] = (x[29]);
  assign t[441] = (x[61]);
  assign t[442] = (x[62]);
  assign t[443] = (x[69]);
  assign t[444] = (x[70]);
  assign t[445] = (x[75]);
  assign t[446] = (x[76]);
  assign t[447] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[448] = (x[106]);
  assign t[449] = (x[37]);
  assign t[44] = ~(t[73] ^ t[74]);
  assign t[450] = (x[45]);
  assign t[451] = (x[86]);
  assign t[452] = (x[87]);
  assign t[453] = (x[51]);
  assign t[454] = (x[59]);
  assign t[455] = (x[67]);
  assign t[456] = (x[73]);
  assign t[457] = (x[107]);
  assign t[458] = (x[108]);
  assign t[459] = (x[84]);
  assign t[45] = ~(t[75] | t[76]);
  assign t[460] = (x[105]);
  assign t[46] = ~(t[47] ^ t[77]);
  assign t[47] = ~(t[78] | t[79]);
  assign t[48] = ~(t[80] ^ t[81]);
  assign t[49] = ~(t[209]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[82] & t[83]);
  assign t[51] = t[84] | t[85];
  assign t[52] = t[210] & t[86];
  assign t[53] = t[87] | t[88];
  assign t[54] = ~(t[213]);
  assign t[55] = ~(t[214]);
  assign t[56] = ~(t[89] | t[90]);
  assign t[57] = ~(t[91] | t[92]);
  assign t[58] = ~(t[215] | t[93]);
  assign t[59] = t[30] ? x[44] : x[43];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[94] & t[95]);
  assign t[61] = ~(t[96] | t[97]);
  assign t[62] = ~(t[216] | t[98]);
  assign t[63] = ~(t[99] | t[100]);
  assign t[64] = ~(t[101] ^ t[102]);
  assign t[65] = ~(t[103] | t[104]);
  assign t[66] = ~(t[217] | t[105]);
  assign t[67] = ~(t[106] ^ t[107]);
  assign t[68] = ~(t[218]);
  assign t[69] = ~(t[219]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[110] | t[111]);
  assign t[72] = ~(t[220] | t[112]);
  assign t[73] = t[30] ? x[66] : x[65];
  assign t[74] = ~(t[113] & t[83]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[221] | t[116]);
  assign t[77] = ~(t[117] ^ t[118]);
  assign t[78] = ~(t[119] | t[120]);
  assign t[79] = ~(t[222] | t[121]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[122] | t[123]);
  assign t[81] = ~(t[124] ^ t[125]);
  assign t[82] = ~(t[86] & t[126]);
  assign t[83] = ~(t[127] & t[128]);
  assign t[84] = ~(t[129] | t[130]);
  assign t[85] = ~(t[129] | t[131]);
  assign t[86] = ~(t[132] | t[207]);
  assign t[87] = ~(x[7] | t[208]);
  assign t[88] = x[7] & t[208];
  assign t[89] = ~(t[223]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[213] | t[214]);
  assign t[91] = ~(t[224]);
  assign t[92] = ~(t[225]);
  assign t[93] = ~(t[133] | t[134]);
  assign t[94] = ~(t[135] | t[136]);
  assign t[95] = ~(t[85] | t[137]);
  assign t[96] = ~(t[226]);
  assign t[97] = ~(t[227]);
  assign t[98] = ~(t[138] | t[139]);
  assign t[99] = ~(t[140] | t[141]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [172:0] x;
 output y;

 wire [667:0] t;
  assign t[0] = t[1] ? t[2] : t[398];
  assign t[100] = t[135] ? x[89] : x[88];
  assign t[101] = ~(t[139] & t[140]);
  assign t[102] = ~(t[422]);
  assign t[103] = ~(t[410] | t[411]);
  assign t[104] = ~(t[423]);
  assign t[105] = ~(t[424]);
  assign t[106] = ~(t[141] | t[142]);
  assign t[107] = ~(t[139] & t[143]);
  assign t[108] = ~(t[425]);
  assign t[109] = ~(t[426]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[144] | t[145]);
  assign t[111] = ~(t[146] | t[147]);
  assign t[112] = ~(t[427] | t[148]);
  assign t[113] = t[149] ? x[102] : x[101];
  assign t[114] = ~(t[150] & t[151]);
  assign t[115] = ~(t[428]);
  assign t[116] = ~(t[429]);
  assign t[117] = ~(t[152] | t[153]);
  assign t[118] = ~(t[154] | t[155]);
  assign t[119] = ~(t[430] | t[156]);
  assign t[11] = ~(x[6]);
  assign t[120] = t[149] ? x[112] : x[111];
  assign t[121] = ~(t[157] & t[143]);
  assign t[122] = ~(t[401]);
  assign t[123] = ~(t[158] & t[159]);
  assign t[124] = ~(t[160] & t[402]);
  assign t[125] = ~(t[81] | t[161]);
  assign t[126] = ~(t[81] | t[162]);
  assign t[127] = ~(x[7] & t[163]);
  assign t[128] = ~(t[402] & t[164]);
  assign t[129] = ~(t[431]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[416] | t[417]);
  assign t[131] = ~(t[157] & t[139]);
  assign t[132] = ~(t[81] | t[165]);
  assign t[133] = ~(t[432]);
  assign t[134] = ~(t[418] | t[419]);
  assign t[135] = ~(t[49]);
  assign t[136] = ~(t[166] | t[167]);
  assign t[137] = ~(t[433]);
  assign t[138] = ~(t[420] | t[421]);
  assign t[139] = ~(t[168] | t[167]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[169] | t[170]);
  assign t[141] = ~(t[434]);
  assign t[142] = ~(t[423] | t[424]);
  assign t[143] = ~(t[171] & t[172]);
  assign t[144] = ~(t[435]);
  assign t[145] = ~(t[425] | t[426]);
  assign t[146] = ~(t[436]);
  assign t[147] = ~(t[437]);
  assign t[148] = ~(t[173] | t[174]);
  assign t[149] = ~(t[49]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[175] | t[176]);
  assign t[151] = ~(t[177] & t[178]);
  assign t[152] = ~(t[438]);
  assign t[153] = ~(t[428] | t[429]);
  assign t[154] = ~(t[439]);
  assign t[155] = ~(t[440]);
  assign t[156] = ~(t[179] | t[180]);
  assign t[157] = ~(t[50] | t[169]);
  assign t[158] = ~(x[7] | t[400]);
  assign t[159] = ~(t[402]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = x[7] & t[400];
  assign t[161] = t[399] ? t[182] : t[181];
  assign t[162] = t[399] ? t[184] : t[183];
  assign t[163] = ~(t[400] | t[402]);
  assign t[164] = ~(x[7] | t[185]);
  assign t[165] = t[399] ? t[123] : t[124];
  assign t[166] = ~(t[122] | t[186]);
  assign t[167] = ~(t[122] | t[187]);
  assign t[168] = ~(t[122] | t[188]);
  assign t[169] = ~(t[189] & t[190]);
  assign t[16] = ~(t[399] & t[400]);
  assign t[170] = ~(t[151] & t[191]);
  assign t[171] = ~(t[400] | t[159]);
  assign t[172] = t[81] & t[399];
  assign t[173] = ~(t[441]);
  assign t[174] = ~(t[436] | t[437]);
  assign t[175] = ~(t[192] & t[143]);
  assign t[176] = t[52] | t[193];
  assign t[177] = t[402] & t[194];
  assign t[178] = t[158] | t[160];
  assign t[179] = ~(t[442]);
  assign t[17] = ~(t[401] & t[402]);
  assign t[180] = ~(t[439] | t[440]);
  assign t[181] = ~(t[164] & t[159]);
  assign t[182] = ~(x[7] & t[171]);
  assign t[183] = ~(t[158] & t[402]);
  assign t[184] = ~(t[160] & t[159]);
  assign t[185] = ~(t[400]);
  assign t[186] = t[399] ? t[123] : t[184];
  assign t[187] = t[399] ? t[181] : t[127];
  assign t[188] = t[399] ? t[184] : t[123];
  assign t[189] = ~(t[166] | t[195]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[122] & t[196]);
  assign t[191] = t[122] | t[197];
  assign t[192] = ~(t[194] & t[198]);
  assign t[193] = ~(t[81] | t[199]);
  assign t[194] = ~(t[122] | t[399]);
  assign t[195] = ~(t[81] | t[200]);
  assign t[196] = ~(t[127] & t[128]);
  assign t[197] = t[399] ? t[127] : t[181];
  assign t[198] = ~(t[128] & t[182]);
  assign t[199] = t[399] ? t[183] : t[184];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[399] ? t[181] : t[182];
  assign t[201] = t[6] ? t[202] : t[443];
  assign t[202] = x[6] ? t[204] : t[203];
  assign t[203] = x[7] ? t[206] : t[205];
  assign t[204] = t[207] ^ x[126];
  assign t[205] = t[208] ^ t[209];
  assign t[206] = ~(t[210] ^ t[211]);
  assign t[207] = x[127] ^ x[128];
  assign t[208] = t[30] ? x[128] : x[127];
  assign t[209] = ~(t[212] ^ t[213]);
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = x[7] ? t[215] : t[214];
  assign t[211] = ~(t[216] ^ t[217]);
  assign t[212] = x[7] ? t[219] : t[218];
  assign t[213] = ~(t[220] ^ t[221]);
  assign t[214] = ~(t[222] & t[223]);
  assign t[215] = t[224] ^ t[225];
  assign t[216] = x[7] ? t[227] : t[226];
  assign t[217] = x[7] ? t[229] : t[228];
  assign t[218] = ~(t[230] & t[231]);
  assign t[219] = t[232] ^ t[233];
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = x[7] ? t[235] : t[234];
  assign t[221] = x[7] ? t[237] : t[236];
  assign t[222] = ~(t[405] & t[54]);
  assign t[223] = ~(t[415] & t[238]);
  assign t[224] = t[30] ? x[130] : x[129];
  assign t[225] = ~(t[239] & t[240]);
  assign t[226] = ~(t[241] & t[242]);
  assign t[227] = t[243] ^ t[234];
  assign t[228] = ~(t[244] & t[245]);
  assign t[229] = t[246] ^ t[228];
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = ~(t[410] & t[67]);
  assign t[231] = ~(t[422] & t[247]);
  assign t[232] = t[30] ? x[132] : x[131];
  assign t[233] = ~(t[248] & t[249]);
  assign t[234] = ~(t[250] & t[251]);
  assign t[235] = t[252] ^ t[253];
  assign t[236] = ~(t[254] & t[255]);
  assign t[237] = t[256] ^ t[257];
  assign t[238] = ~(t[406] & t[53]);
  assign t[239] = ~(t[416] & t[88]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = ~(t[431] & t[258]);
  assign t[241] = ~(t[420] & t[98]);
  assign t[242] = ~(t[433] & t[259]);
  assign t[243] = t[135] ? x[134] : x[133];
  assign t[244] = ~(t[418] & t[93]);
  assign t[245] = ~(t[432] & t[260]);
  assign t[246] = t[135] ? x[136] : x[135];
  assign t[247] = ~(t[411] & t[66]);
  assign t[248] = ~(t[423] & t[105]);
  assign t[249] = ~(t[434] & t[261]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = ~(t[428] & t[116]);
  assign t[251] = ~(t[438] & t[262]);
  assign t[252] = t[149] ? x[138] : x[137];
  assign t[253] = ~(t[263] & t[264]);
  assign t[254] = ~(t[425] & t[109]);
  assign t[255] = ~(t[435] & t[265]);
  assign t[256] = t[149] ? x[140] : x[139];
  assign t[257] = ~(t[266] & t[267]);
  assign t[258] = ~(t[417] & t[87]);
  assign t[259] = ~(t[421] & t[97]);
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = ~(t[419] & t[92]);
  assign t[261] = ~(t[424] & t[104]);
  assign t[262] = ~(t[429] & t[115]);
  assign t[263] = ~(t[439] & t[155]);
  assign t[264] = ~(t[442] & t[268]);
  assign t[265] = ~(t[426] & t[108]);
  assign t[266] = ~(t[436] & t[147]);
  assign t[267] = ~(t[441] & t[269]);
  assign t[268] = ~(t[440] & t[154]);
  assign t[269] = ~(t[437] & t[146]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[6] ? t[271] : t[444];
  assign t[271] = x[6] ? t[273] : t[272];
  assign t[272] = x[7] ? t[275] : t[274];
  assign t[273] = t[276] ^ x[142];
  assign t[274] = t[277] ^ t[278];
  assign t[275] = ~(t[279] ^ t[280]);
  assign t[276] = x[143] ^ x[144];
  assign t[277] = t[30] ? x[144] : x[143];
  assign t[278] = ~(t[281] ^ t[282]);
  assign t[279] = x[7] ? t[284] : t[283];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = ~(t[285] ^ t[286]);
  assign t[281] = x[7] ? t[288] : t[287];
  assign t[282] = ~(t[289] ^ t[290]);
  assign t[283] = ~(t[291] & t[292]);
  assign t[284] = t[293] ^ t[294];
  assign t[285] = x[7] ? t[296] : t[295];
  assign t[286] = x[7] ? t[298] : t[297];
  assign t[287] = ~(t[299] & t[300]);
  assign t[288] = t[301] ^ t[302];
  assign t[289] = x[7] ? t[304] : t[303];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = x[7] ? t[306] : t[305];
  assign t[291] = ~(t[54] & t[85]);
  assign t[292] = ~(t[307] & t[403]);
  assign t[293] = t[30] ? x[146] : x[145];
  assign t[294] = ~(t[308] & t[309]);
  assign t[295] = ~(t[310] & t[311]);
  assign t[296] = t[312] ^ t[295];
  assign t[297] = ~(t[313] & t[314]);
  assign t[298] = t[315] ^ t[303];
  assign t[299] = ~(t[67] & t[102]);
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = ~(t[316] & t[404]);
  assign t[301] = t[30] ? x[148] : x[147];
  assign t[302] = ~(t[317] & t[318]);
  assign t[303] = ~(t[319] & t[320]);
  assign t[304] = t[321] ^ t[322];
  assign t[305] = ~(t[323] & t[324]);
  assign t[306] = t[325] ^ t[326];
  assign t[307] = ~(t[327] & t[53]);
  assign t[308] = ~(t[88] & t[129]);
  assign t[309] = ~(t[328] & t[407]);
  assign t[30] = ~(t[49]);
  assign t[310] = ~(t[93] & t[133]);
  assign t[311] = ~(t[329] & t[408]);
  assign t[312] = t[135] ? x[150] : x[149];
  assign t[313] = ~(t[98] & t[137]);
  assign t[314] = ~(t[330] & t[409]);
  assign t[315] = t[135] ? x[152] : x[151];
  assign t[316] = ~(t[331] & t[66]);
  assign t[317] = ~(t[105] & t[141]);
  assign t[318] = ~(t[332] & t[412]);
  assign t[319] = ~(t[116] & t[152]);
  assign t[31] = ~(t[50]);
  assign t[320] = ~(t[333] & t[414]);
  assign t[321] = t[149] ? x[154] : x[153];
  assign t[322] = ~(t[334] & t[335]);
  assign t[323] = ~(t[109] & t[144]);
  assign t[324] = ~(t[336] & t[413]);
  assign t[325] = t[149] ? x[156] : x[155];
  assign t[326] = ~(t[337] & t[338]);
  assign t[327] = ~(t[415] & t[406]);
  assign t[328] = ~(t[339] & t[87]);
  assign t[329] = ~(t[340] & t[92]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = ~(t[341] & t[97]);
  assign t[331] = ~(t[422] & t[411]);
  assign t[332] = ~(t[342] & t[104]);
  assign t[333] = ~(t[343] & t[115]);
  assign t[334] = ~(t[155] & t[179]);
  assign t[335] = ~(t[344] & t[430]);
  assign t[336] = ~(t[345] & t[108]);
  assign t[337] = ~(t[147] & t[173]);
  assign t[338] = ~(t[346] & t[427]);
  assign t[339] = ~(t[431] & t[417]);
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = ~(t[432] & t[419]);
  assign t[341] = ~(t[433] & t[421]);
  assign t[342] = ~(t[434] & t[424]);
  assign t[343] = ~(t[438] & t[429]);
  assign t[344] = ~(t[347] & t[154]);
  assign t[345] = ~(t[435] & t[426]);
  assign t[346] = ~(t[348] & t[146]);
  assign t[347] = ~(t[442] & t[440]);
  assign t[348] = ~(t[441] & t[437]);
  assign t[349] = t[1] ? t[350] : t[445];
  assign t[34] = ~(t[403] | t[55]);
  assign t[350] = x[6] ? t[352] : t[351];
  assign t[351] = x[7] ? t[354] : t[353];
  assign t[352] = t[355] ^ x[158];
  assign t[353] = t[356] ^ t[357];
  assign t[354] = ~(t[358] ^ t[359]);
  assign t[355] = x[159] ^ x[160];
  assign t[356] = t[30] ? x[160] : x[159];
  assign t[357] = ~(t[360] ^ t[361]);
  assign t[358] = x[7] ? t[363] : t[362];
  assign t[359] = ~(t[364] ^ t[365]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = x[7] ? t[367] : t[366];
  assign t[361] = ~(t[368] ^ t[369]);
  assign t[362] = ~(t[291] & t[370]);
  assign t[363] = t[371] ^ t[372];
  assign t[364] = x[7] ? t[374] : t[373];
  assign t[365] = x[7] ? t[376] : t[375];
  assign t[366] = ~(t[299] & t[377]);
  assign t[367] = t[378] ^ t[379];
  assign t[368] = x[7] ? t[381] : t[380];
  assign t[369] = x[7] ? t[383] : t[382];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[33] | t[403];
  assign t[371] = t[30] ? x[162] : x[161];
  assign t[372] = ~(t[308] & t[384]);
  assign t[373] = ~(t[310] & t[385]);
  assign t[374] = t[386] ^ t[373];
  assign t[375] = ~(t[313] & t[387]);
  assign t[376] = t[388] ^ t[380];
  assign t[377] = t[41] | t[404];
  assign t[378] = t[30] ? x[164] : x[163];
  assign t[379] = ~(t[317] & t[389]);
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = ~(t[319] & t[390]);
  assign t[381] = t[391] ^ t[392];
  assign t[382] = ~(t[323] & t[393]);
  assign t[383] = t[394] ^ t[395];
  assign t[384] = t[56] | t[407];
  assign t[385] = t[60] | t[408];
  assign t[386] = t[135] ? x[166] : x[165];
  assign t[387] = t[63] | t[409];
  assign t[388] = t[135] ? x[168] : x[167];
  assign t[389] = t[69] | t[412];
  assign t[38] = ~(t[37] ^ t[62]);
  assign t[390] = t[77] | t[414];
  assign t[391] = t[149] ? x[170] : x[169];
  assign t[392] = ~(t[334] & t[396]);
  assign t[393] = t[73] | t[413];
  assign t[394] = t[149] ? x[172] : x[171];
  assign t[395] = ~(t[337] & t[397]);
  assign t[396] = t[118] | t[430];
  assign t[397] = t[111] | t[427];
  assign t[398] = (t[446]);
  assign t[399] = (t[447]);
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (t[448]);
  assign t[401] = (t[449]);
  assign t[402] = (t[450]);
  assign t[403] = (t[451]);
  assign t[404] = (t[452]);
  assign t[405] = (t[453]);
  assign t[406] = (t[454]);
  assign t[407] = (t[455]);
  assign t[408] = (t[456]);
  assign t[409] = (t[457]);
  assign t[40] = ~(t[47] ^ t[65]);
  assign t[410] = (t[458]);
  assign t[411] = (t[459]);
  assign t[412] = (t[460]);
  assign t[413] = (t[461]);
  assign t[414] = (t[462]);
  assign t[415] = (t[463]);
  assign t[416] = (t[464]);
  assign t[417] = (t[465]);
  assign t[418] = (t[466]);
  assign t[419] = (t[467]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (t[468]);
  assign t[421] = (t[469]);
  assign t[422] = (t[470]);
  assign t[423] = (t[471]);
  assign t[424] = (t[472]);
  assign t[425] = (t[473]);
  assign t[426] = (t[474]);
  assign t[427] = (t[475]);
  assign t[428] = (t[476]);
  assign t[429] = (t[477]);
  assign t[42] = ~(t[404] | t[68]);
  assign t[430] = (t[478]);
  assign t[431] = (t[479]);
  assign t[432] = (t[480]);
  assign t[433] = (t[481]);
  assign t[434] = (t[482]);
  assign t[435] = (t[483]);
  assign t[436] = (t[484]);
  assign t[437] = (t[485]);
  assign t[438] = (t[486]);
  assign t[439] = (t[487]);
  assign t[43] = ~(t[69] | t[70]);
  assign t[440] = (t[488]);
  assign t[441] = (t[489]);
  assign t[442] = (t[490]);
  assign t[443] = (t[491]);
  assign t[444] = (t[492]);
  assign t[445] = (t[493]);
  assign t[446] = t[494] ^ x[5];
  assign t[447] = t[495] ^ x[13];
  assign t[448] = t[496] ^ x[16];
  assign t[449] = t[497] ^ x[19];
  assign t[44] = ~(t[71] ^ t[72]);
  assign t[450] = t[498] ^ x[22];
  assign t[451] = t[499] ^ x[28];
  assign t[452] = t[500] ^ x[34];
  assign t[453] = t[501] ^ x[35];
  assign t[454] = t[502] ^ x[36];
  assign t[455] = t[503] ^ x[42];
  assign t[456] = t[504] ^ x[50];
  assign t[457] = t[505] ^ x[56];
  assign t[458] = t[506] ^ x[57];
  assign t[459] = t[507] ^ x[58];
  assign t[45] = ~(t[73] | t[74]);
  assign t[460] = t[508] ^ x[64];
  assign t[461] = t[509] ^ x[72];
  assign t[462] = t[510] ^ x[78];
  assign t[463] = t[511] ^ x[79];
  assign t[464] = t[512] ^ x[80];
  assign t[465] = t[513] ^ x[81];
  assign t[466] = t[514] ^ x[82];
  assign t[467] = t[515] ^ x[83];
  assign t[468] = t[516] ^ x[86];
  assign t[469] = t[517] ^ x[87];
  assign t[46] = ~(t[75] ^ t[76]);
  assign t[470] = t[518] ^ x[90];
  assign t[471] = t[519] ^ x[91];
  assign t[472] = t[520] ^ x[92];
  assign t[473] = t[521] ^ x[93];
  assign t[474] = t[522] ^ x[94];
  assign t[475] = t[523] ^ x[100];
  assign t[476] = t[524] ^ x[103];
  assign t[477] = t[525] ^ x[104];
  assign t[478] = t[526] ^ x[110];
  assign t[479] = t[527] ^ x[113];
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = t[528] ^ x[114];
  assign t[481] = t[529] ^ x[115];
  assign t[482] = t[530] ^ x[116];
  assign t[483] = t[531] ^ x[117];
  assign t[484] = t[532] ^ x[118];
  assign t[485] = t[533] ^ x[119];
  assign t[486] = t[534] ^ x[120];
  assign t[487] = t[535] ^ x[121];
  assign t[488] = t[536] ^ x[122];
  assign t[489] = t[537] ^ x[123];
  assign t[48] = ~(t[79] ^ t[80]);
  assign t[490] = t[538] ^ x[124];
  assign t[491] = t[539] ^ x[125];
  assign t[492] = t[540] ^ x[141];
  assign t[493] = t[541] ^ x[157];
  assign t[494] = (~t[542] & t[543]);
  assign t[495] = (~t[544] & t[545]);
  assign t[496] = (~t[546] & t[547]);
  assign t[497] = (~t[548] & t[549]);
  assign t[498] = (~t[550] & t[551]);
  assign t[499] = (~t[552] & t[553]);
  assign t[49] = ~(t[401]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[554] & t[555]);
  assign t[501] = (~t[552] & t[556]);
  assign t[502] = (~t[552] & t[557]);
  assign t[503] = (~t[558] & t[559]);
  assign t[504] = (~t[560] & t[561]);
  assign t[505] = (~t[562] & t[563]);
  assign t[506] = (~t[554] & t[564]);
  assign t[507] = (~t[554] & t[565]);
  assign t[508] = (~t[566] & t[567]);
  assign t[509] = (~t[568] & t[569]);
  assign t[50] = ~(t[81] | t[82]);
  assign t[510] = (~t[570] & t[571]);
  assign t[511] = (~t[552] & t[572]);
  assign t[512] = (~t[558] & t[573]);
  assign t[513] = (~t[558] & t[574]);
  assign t[514] = (~t[560] & t[575]);
  assign t[515] = (~t[560] & t[576]);
  assign t[516] = (~t[562] & t[577]);
  assign t[517] = (~t[562] & t[578]);
  assign t[518] = (~t[554] & t[579]);
  assign t[519] = (~t[566] & t[580]);
  assign t[51] = ~(t[83]);
  assign t[520] = (~t[566] & t[581]);
  assign t[521] = (~t[568] & t[582]);
  assign t[522] = (~t[568] & t[583]);
  assign t[523] = (~t[584] & t[585]);
  assign t[524] = (~t[570] & t[586]);
  assign t[525] = (~t[570] & t[587]);
  assign t[526] = (~t[588] & t[589]);
  assign t[527] = (~t[558] & t[590]);
  assign t[528] = (~t[560] & t[591]);
  assign t[529] = (~t[562] & t[592]);
  assign t[52] = ~(t[81] | t[84]);
  assign t[530] = (~t[566] & t[593]);
  assign t[531] = (~t[568] & t[594]);
  assign t[532] = (~t[584] & t[595]);
  assign t[533] = (~t[584] & t[596]);
  assign t[534] = (~t[570] & t[597]);
  assign t[535] = (~t[588] & t[598]);
  assign t[536] = (~t[588] & t[599]);
  assign t[537] = (~t[584] & t[600]);
  assign t[538] = (~t[588] & t[601]);
  assign t[539] = (~t[542] & t[602]);
  assign t[53] = ~(t[405]);
  assign t[540] = (~t[542] & t[603]);
  assign t[541] = (~t[542] & t[604]);
  assign t[542] = t[605] ^ x[4];
  assign t[543] = t[606] ^ x[5];
  assign t[544] = t[607] ^ x[12];
  assign t[545] = t[608] ^ x[13];
  assign t[546] = t[609] ^ x[15];
  assign t[547] = t[610] ^ x[16];
  assign t[548] = t[611] ^ x[18];
  assign t[549] = t[612] ^ x[19];
  assign t[54] = ~(t[406]);
  assign t[550] = t[613] ^ x[21];
  assign t[551] = t[614] ^ x[22];
  assign t[552] = t[615] ^ x[27];
  assign t[553] = t[616] ^ x[28];
  assign t[554] = t[617] ^ x[33];
  assign t[555] = t[618] ^ x[34];
  assign t[556] = t[619] ^ x[35];
  assign t[557] = t[620] ^ x[36];
  assign t[558] = t[621] ^ x[41];
  assign t[559] = t[622] ^ x[42];
  assign t[55] = ~(t[85] | t[86]);
  assign t[560] = t[623] ^ x[49];
  assign t[561] = t[624] ^ x[50];
  assign t[562] = t[625] ^ x[55];
  assign t[563] = t[626] ^ x[56];
  assign t[564] = t[627] ^ x[57];
  assign t[565] = t[628] ^ x[58];
  assign t[566] = t[629] ^ x[63];
  assign t[567] = t[630] ^ x[64];
  assign t[568] = t[631] ^ x[71];
  assign t[569] = t[632] ^ x[72];
  assign t[56] = ~(t[87] | t[88]);
  assign t[570] = t[633] ^ x[77];
  assign t[571] = t[634] ^ x[78];
  assign t[572] = t[635] ^ x[79];
  assign t[573] = t[636] ^ x[80];
  assign t[574] = t[637] ^ x[81];
  assign t[575] = t[638] ^ x[82];
  assign t[576] = t[639] ^ x[83];
  assign t[577] = t[640] ^ x[86];
  assign t[578] = t[641] ^ x[87];
  assign t[579] = t[642] ^ x[90];
  assign t[57] = ~(t[407] | t[89]);
  assign t[580] = t[643] ^ x[91];
  assign t[581] = t[644] ^ x[92];
  assign t[582] = t[645] ^ x[93];
  assign t[583] = t[646] ^ x[94];
  assign t[584] = t[647] ^ x[99];
  assign t[585] = t[648] ^ x[100];
  assign t[586] = t[649] ^ x[103];
  assign t[587] = t[650] ^ x[104];
  assign t[588] = t[651] ^ x[109];
  assign t[589] = t[652] ^ x[110];
  assign t[58] = t[30] ? x[44] : x[43];
  assign t[590] = t[653] ^ x[113];
  assign t[591] = t[654] ^ x[114];
  assign t[592] = t[655] ^ x[115];
  assign t[593] = t[656] ^ x[116];
  assign t[594] = t[657] ^ x[117];
  assign t[595] = t[658] ^ x[118];
  assign t[596] = t[659] ^ x[119];
  assign t[597] = t[660] ^ x[120];
  assign t[598] = t[661] ^ x[121];
  assign t[599] = t[662] ^ x[122];
  assign t[59] = ~(t[90] & t[91]);
  assign t[5] = t[9] ^ x[8];
  assign t[600] = t[663] ^ x[123];
  assign t[601] = t[664] ^ x[124];
  assign t[602] = t[665] ^ x[125];
  assign t[603] = t[666] ^ x[141];
  assign t[604] = t[667] ^ x[157];
  assign t[605] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[606] = (x[0]);
  assign t[607] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[608] = (x[11]);
  assign t[609] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[60] = ~(t[92] | t[93]);
  assign t[610] = (x[14]);
  assign t[611] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[612] = (x[17]);
  assign t[613] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[614] = (x[20]);
  assign t[615] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[616] = (x[24]);
  assign t[617] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[618] = (x[30]);
  assign t[619] = (x[25]);
  assign t[61] = ~(t[408] | t[94]);
  assign t[620] = (x[26]);
  assign t[621] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[622] = (x[38]);
  assign t[623] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[624] = (x[46]);
  assign t[625] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[626] = (x[52]);
  assign t[627] = (x[31]);
  assign t[628] = (x[32]);
  assign t[629] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[62] = ~(t[95] ^ t[96]);
  assign t[630] = (x[60]);
  assign t[631] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[632] = (x[68]);
  assign t[633] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[634] = (x[74]);
  assign t[635] = (x[23]);
  assign t[636] = (x[39]);
  assign t[637] = (x[40]);
  assign t[638] = (x[47]);
  assign t[639] = (x[48]);
  assign t[63] = ~(t[97] | t[98]);
  assign t[640] = (x[53]);
  assign t[641] = (x[54]);
  assign t[642] = (x[29]);
  assign t[643] = (x[61]);
  assign t[644] = (x[62]);
  assign t[645] = (x[69]);
  assign t[646] = (x[70]);
  assign t[647] = (x[95] & ~x[96] & ~x[97] & ~x[98]) | (~x[95] & x[96] & ~x[97] & ~x[98]) | (~x[95] & ~x[96] & x[97] & ~x[98]) | (~x[95] & ~x[96] & ~x[97] & x[98]) | (x[95] & x[96] & x[97] & ~x[98]) | (x[95] & x[96] & ~x[97] & x[98]) | (x[95] & ~x[96] & x[97] & x[98]) | (~x[95] & x[96] & x[97] & x[98]);
  assign t[648] = (x[96]);
  assign t[649] = (x[75]);
  assign t[64] = ~(t[409] | t[99]);
  assign t[650] = (x[76]);
  assign t[651] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[652] = (x[106]);
  assign t[653] = (x[37]);
  assign t[654] = (x[45]);
  assign t[655] = (x[51]);
  assign t[656] = (x[59]);
  assign t[657] = (x[67]);
  assign t[658] = (x[97]);
  assign t[659] = (x[98]);
  assign t[65] = ~(t[100] ^ t[101]);
  assign t[660] = (x[73]);
  assign t[661] = (x[107]);
  assign t[662] = (x[108]);
  assign t[663] = (x[95]);
  assign t[664] = (x[105]);
  assign t[665] = (x[1]);
  assign t[666] = (x[2]);
  assign t[667] = (x[3]);
  assign t[66] = ~(t[410]);
  assign t[67] = ~(t[411]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[104] | t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[412] | t[106]);
  assign t[71] = t[30] ? x[66] : x[65];
  assign t[72] = t[107] | t[52];
  assign t[73] = ~(t[108] | t[109]);
  assign t[74] = ~(t[413] | t[110]);
  assign t[75] = ~(t[111] | t[112]);
  assign t[76] = ~(t[113] ^ t[114]);
  assign t[77] = ~(t[115] | t[116]);
  assign t[78] = ~(t[414] | t[117]);
  assign t[79] = ~(t[118] | t[119]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[120] ^ t[121]);
  assign t[81] = ~(t[122]);
  assign t[82] = t[399] ? t[124] : t[123];
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = t[399] ? t[128] : t[127];
  assign t[85] = ~(t[415]);
  assign t[86] = ~(t[405] | t[406]);
  assign t[87] = ~(t[416]);
  assign t[88] = ~(t[417]);
  assign t[89] = ~(t[129] | t[130]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125] | t[131]);
  assign t[91] = ~(t[132]);
  assign t[92] = ~(t[418]);
  assign t[93] = ~(t[419]);
  assign t[94] = ~(t[133] | t[134]);
  assign t[95] = t[135] ? x[85] : x[84];
  assign t[96] = ~(t[136] & t[32]);
  assign t[97] = ~(t[420]);
  assign t[98] = ~(t[421]);
  assign t[99] = ~(t[137] | t[138]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[201] & ~t[270] & ~t[349]) | (~t[0] & t[201] & ~t[270] & ~t[349]) | (~t[0] & ~t[201] & t[270] & ~t[349]) | (~t[0] & ~t[201] & ~t[270] & t[349]) | (t[0] & t[201] & t[270] & ~t[349]) | (t[0] & t[201] & ~t[270] & t[349]) | (t[0] & ~t[201] & t[270] & t[349]) | (~t[0] & t[201] & t[270] & t[349]);
endmodule

module R2ind161(x, y);
 input [124:0] x;
 output y;

 wire [364:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[147]);
  assign t[101] = ~(t[148]);
  assign t[102] = ~(t[149]);
  assign t[103] = ~(t[108] | t[101]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[5];
  assign t[156] = t[201] ^ x[13];
  assign t[157] = t[202] ^ x[16];
  assign t[158] = t[203] ^ x[19];
  assign t[159] = t[204] ^ x[22];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[28];
  assign t[161] = t[206] ^ x[36];
  assign t[162] = t[207] ^ x[39];
  assign t[163] = t[208] ^ x[40];
  assign t[164] = t[209] ^ x[46];
  assign t[165] = t[210] ^ x[52];
  assign t[166] = t[211] ^ x[60];
  assign t[167] = t[212] ^ x[63];
  assign t[168] = t[213] ^ x[64];
  assign t[169] = t[214] ^ x[70];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[76];
  assign t[171] = t[216] ^ x[84];
  assign t[172] = t[217] ^ x[87];
  assign t[173] = t[218] ^ x[88];
  assign t[174] = t[219] ^ x[89];
  assign t[175] = t[220] ^ x[90];
  assign t[176] = t[221] ^ x[91];
  assign t[177] = t[222] ^ x[92];
  assign t[178] = t[223] ^ x[93];
  assign t[179] = t[224] ^ x[94];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[95];
  assign t[181] = t[226] ^ x[96];
  assign t[182] = t[227] ^ x[97];
  assign t[183] = t[228] ^ x[98];
  assign t[184] = t[229] ^ x[104];
  assign t[185] = t[230] ^ x[105];
  assign t[186] = t[231] ^ x[106];
  assign t[187] = t[232] ^ x[112];
  assign t[188] = t[233] ^ x[113];
  assign t[189] = t[234] ^ x[114];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[115];
  assign t[191] = t[236] ^ x[116];
  assign t[192] = t[237] ^ x[117];
  assign t[193] = t[238] ^ x[118];
  assign t[194] = t[239] ^ x[119];
  assign t[195] = t[240] ^ x[120];
  assign t[196] = t[241] ^ x[121];
  assign t[197] = t[242] ^ x[122];
  assign t[198] = t[243] ^ x[123];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[245] & t[246]);
  assign t[201] = (~t[247] & t[248]);
  assign t[202] = (~t[249] & t[250]);
  assign t[203] = (~t[251] & t[252]);
  assign t[204] = (~t[253] & t[254]);
  assign t[205] = (~t[255] & t[256]);
  assign t[206] = (~t[257] & t[258]);
  assign t[207] = (~t[255] & t[259]);
  assign t[208] = (~t[255] & t[260]);
  assign t[209] = (~t[261] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[263] & t[264]);
  assign t[211] = (~t[265] & t[266]);
  assign t[212] = (~t[257] & t[267]);
  assign t[213] = (~t[257] & t[268]);
  assign t[214] = (~t[269] & t[270]);
  assign t[215] = (~t[271] & t[272]);
  assign t[216] = (~t[273] & t[274]);
  assign t[217] = (~t[255] & t[275]);
  assign t[218] = (~t[261] & t[276]);
  assign t[219] = (~t[261] & t[277]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[263] & t[278]);
  assign t[221] = (~t[263] & t[279]);
  assign t[222] = (~t[265] & t[280]);
  assign t[223] = (~t[265] & t[281]);
  assign t[224] = (~t[257] & t[282]);
  assign t[225] = (~t[269] & t[283]);
  assign t[226] = (~t[269] & t[284]);
  assign t[227] = (~t[271] & t[285]);
  assign t[228] = (~t[271] & t[286]);
  assign t[229] = (~t[287] & t[288]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[273] & t[289]);
  assign t[231] = (~t[273] & t[290]);
  assign t[232] = (~t[291] & t[292]);
  assign t[233] = (~t[261] & t[293]);
  assign t[234] = (~t[263] & t[294]);
  assign t[235] = (~t[265] & t[295]);
  assign t[236] = (~t[269] & t[296]);
  assign t[237] = (~t[271] & t[297]);
  assign t[238] = (~t[287] & t[298]);
  assign t[239] = (~t[287] & t[299]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[273] & t[300]);
  assign t[241] = (~t[291] & t[301]);
  assign t[242] = (~t[291] & t[302]);
  assign t[243] = (~t[287] & t[303]);
  assign t[244] = (~t[291] & t[304]);
  assign t[245] = t[305] ^ x[4];
  assign t[246] = t[306] ^ x[5];
  assign t[247] = t[307] ^ x[12];
  assign t[248] = t[308] ^ x[13];
  assign t[249] = t[309] ^ x[15];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[310] ^ x[16];
  assign t[251] = t[311] ^ x[18];
  assign t[252] = t[312] ^ x[19];
  assign t[253] = t[313] ^ x[21];
  assign t[254] = t[314] ^ x[22];
  assign t[255] = t[315] ^ x[27];
  assign t[256] = t[316] ^ x[28];
  assign t[257] = t[317] ^ x[35];
  assign t[258] = t[318] ^ x[36];
  assign t[259] = t[319] ^ x[39];
  assign t[25] = ~(t[113]);
  assign t[260] = t[320] ^ x[40];
  assign t[261] = t[321] ^ x[45];
  assign t[262] = t[322] ^ x[46];
  assign t[263] = t[323] ^ x[51];
  assign t[264] = t[324] ^ x[52];
  assign t[265] = t[325] ^ x[59];
  assign t[266] = t[326] ^ x[60];
  assign t[267] = t[327] ^ x[63];
  assign t[268] = t[328] ^ x[64];
  assign t[269] = t[329] ^ x[69];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[70];
  assign t[271] = t[331] ^ x[75];
  assign t[272] = t[332] ^ x[76];
  assign t[273] = t[333] ^ x[83];
  assign t[274] = t[334] ^ x[84];
  assign t[275] = t[335] ^ x[87];
  assign t[276] = t[336] ^ x[88];
  assign t[277] = t[337] ^ x[89];
  assign t[278] = t[338] ^ x[90];
  assign t[279] = t[339] ^ x[91];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[92];
  assign t[281] = t[341] ^ x[93];
  assign t[282] = t[342] ^ x[94];
  assign t[283] = t[343] ^ x[95];
  assign t[284] = t[344] ^ x[96];
  assign t[285] = t[345] ^ x[97];
  assign t[286] = t[346] ^ x[98];
  assign t[287] = t[347] ^ x[103];
  assign t[288] = t[348] ^ x[104];
  assign t[289] = t[349] ^ x[105];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[106];
  assign t[291] = t[351] ^ x[111];
  assign t[292] = t[352] ^ x[112];
  assign t[293] = t[353] ^ x[113];
  assign t[294] = t[354] ^ x[114];
  assign t[295] = t[355] ^ x[115];
  assign t[296] = t[356] ^ x[116];
  assign t[297] = t[357] ^ x[117];
  assign t[298] = t[358] ^ x[118];
  assign t[299] = t[359] ^ x[119];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[120];
  assign t[301] = t[361] ^ x[121];
  assign t[302] = t[362] ^ x[122];
  assign t[303] = t[363] ^ x[123];
  assign t[304] = t[364] ^ x[124];
  assign t[305] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[306] = (x[3]);
  assign t[307] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[308] = (x[11]);
  assign t[309] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = (x[14]);
  assign t[311] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[312] = (x[17]);
  assign t[313] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[314] = (x[20]);
  assign t[315] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[316] = (x[24]);
  assign t[317] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[318] = (x[32]);
  assign t[319] = (x[26]);
  assign t[31] = t[48] | t[115];
  assign t[320] = (x[23]);
  assign t[321] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[322] = (x[42]);
  assign t[323] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[324] = (x[48]);
  assign t[325] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[326] = (x[56]);
  assign t[327] = (x[34]);
  assign t[328] = (x[31]);
  assign t[329] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[32] = t[18] ? x[30] : x[29];
  assign t[330] = (x[66]);
  assign t[331] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[332] = (x[72]);
  assign t[333] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[334] = (x[80]);
  assign t[335] = (x[25]);
  assign t[336] = (x[44]);
  assign t[337] = (x[41]);
  assign t[338] = (x[50]);
  assign t[339] = (x[47]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[58]);
  assign t[341] = (x[55]);
  assign t[342] = (x[33]);
  assign t[343] = (x[68]);
  assign t[344] = (x[65]);
  assign t[345] = (x[74]);
  assign t[346] = (x[71]);
  assign t[347] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[348] = (x[100]);
  assign t[349] = (x[82]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[350] = (x[79]);
  assign t[351] = (x[107] & ~x[108] & ~x[109] & ~x[110]) | (~x[107] & x[108] & ~x[109] & ~x[110]) | (~x[107] & ~x[108] & x[109] & ~x[110]) | (~x[107] & ~x[108] & ~x[109] & x[110]) | (x[107] & x[108] & x[109] & ~x[110]) | (x[107] & x[108] & ~x[109] & x[110]) | (x[107] & ~x[108] & x[109] & x[110]) | (~x[107] & x[108] & x[109] & x[110]);
  assign t[352] = (x[108]);
  assign t[353] = (x[43]);
  assign t[354] = (x[49]);
  assign t[355] = (x[57]);
  assign t[356] = (x[67]);
  assign t[357] = (x[73]);
  assign t[358] = (x[102]);
  assign t[359] = (x[99]);
  assign t[35] = t[53] ^ t[34];
  assign t[360] = (x[81]);
  assign t[361] = (x[110]);
  assign t[362] = (x[107]);
  assign t[363] = (x[101]);
  assign t[364] = (x[109]);
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[42];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = t[59] | t[116];
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[38] : x[37];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[66] & t[67]);
  assign t[45] = t[68] ^ t[69];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[70] | t[46]);
  assign t[49] = ~(t[71] & t[72]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[73] | t[119];
  assign t[51] = ~(t[74] & t[75]);
  assign t[52] = t[76] | t[120];
  assign t[53] = t[77] ? x[54] : x[53];
  assign t[54] = ~(t[78] & t[79]);
  assign t[55] = t[80] | t[121];
  assign t[56] = t[77] ? x[62] : x[61];
  assign t[57] = ~(t[122]);
  assign t[58] = ~(t[123]);
  assign t[59] = ~(t[81] | t[57]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = t[84] | t[124];
  assign t[62] = ~(t[85] & t[86]);
  assign t[63] = t[87] | t[125];
  assign t[64] = t[88] ? x[78] : x[77];
  assign t[65] = ~(t[89] & t[90]);
  assign t[66] = ~(t[91] & t[92]);
  assign t[67] = t[93] | t[126];
  assign t[68] = t[88] ? x[86] : x[85];
  assign t[69] = ~(t[94] & t[95]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[127]);
  assign t[71] = ~(t[128]);
  assign t[72] = ~(t[129]);
  assign t[73] = ~(t[96] | t[71]);
  assign t[74] = ~(t[130]);
  assign t[75] = ~(t[131]);
  assign t[76] = ~(t[97] | t[74]);
  assign t[77] = ~(t[25]);
  assign t[78] = ~(t[132]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[98] | t[78]);
  assign t[81] = ~(t[134]);
  assign t[82] = ~(t[135]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[99] | t[82]);
  assign t[85] = ~(t[137]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[100] | t[85]);
  assign t[88] = ~(t[25]);
  assign t[89] = ~(t[101] & t[102]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = t[103] | t[139];
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [124:0] x;
 output y;

 wire [372:0] t;
  assign t[0] = t[1] ? t[2] : t[118];
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[153]);
  assign t[102] = ~(t[144] & t[143]);
  assign t[103] = ~(t[154]);
  assign t[104] = ~(t[146] & t[145]);
  assign t[105] = ~(t[155]);
  assign t[106] = ~(t[156]);
  assign t[107] = ~(t[157]);
  assign t[108] = ~(t[114] & t[115]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = ~(t[158]);
  assign t[111] = ~(t[159]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[116] & t[117]);
  assign t[114] = ~(t[157] & t[156]);
  assign t[115] = ~(t[161]);
  assign t[116] = ~(t[160] & t[159]);
  assign t[117] = ~(t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[16] ? x[22] : x[21];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[20] : t[19];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = t[208] ^ x[5];
  assign t[164] = t[209] ^ x[11];
  assign t[165] = t[210] ^ x[14];
  assign t[166] = t[211] ^ x[17];
  assign t[167] = t[212] ^ x[20];
  assign t[168] = t[213] ^ x[28];
  assign t[169] = t[214] ^ x[36];
  assign t[16] = ~(t[23]);
  assign t[170] = t[215] ^ x[39];
  assign t[171] = t[216] ^ x[40];
  assign t[172] = t[217] ^ x[46];
  assign t[173] = t[218] ^ x[52];
  assign t[174] = t[219] ^ x[60];
  assign t[175] = t[220] ^ x[63];
  assign t[176] = t[221] ^ x[64];
  assign t[177] = t[222] ^ x[70];
  assign t[178] = t[223] ^ x[76];
  assign t[179] = t[224] ^ x[84];
  assign t[17] = x[7] ? t[25] : t[24];
  assign t[180] = t[225] ^ x[87];
  assign t[181] = t[226] ^ x[88];
  assign t[182] = t[227] ^ x[89];
  assign t[183] = t[228] ^ x[90];
  assign t[184] = t[229] ^ x[91];
  assign t[185] = t[230] ^ x[92];
  assign t[186] = t[231] ^ x[93];
  assign t[187] = t[232] ^ x[94];
  assign t[188] = t[233] ^ x[95];
  assign t[189] = t[234] ^ x[96];
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = t[235] ^ x[97];
  assign t[191] = t[236] ^ x[98];
  assign t[192] = t[237] ^ x[104];
  assign t[193] = t[238] ^ x[105];
  assign t[194] = t[239] ^ x[106];
  assign t[195] = t[240] ^ x[112];
  assign t[196] = t[241] ^ x[113];
  assign t[197] = t[242] ^ x[114];
  assign t[198] = t[243] ^ x[115];
  assign t[199] = t[244] ^ x[116];
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[245] ^ x[117];
  assign t[201] = t[246] ^ x[118];
  assign t[202] = t[247] ^ x[119];
  assign t[203] = t[248] ^ x[120];
  assign t[204] = t[249] ^ x[121];
  assign t[205] = t[250] ^ x[122];
  assign t[206] = t[251] ^ x[123];
  assign t[207] = t[252] ^ x[124];
  assign t[208] = (~t[253] & t[254]);
  assign t[209] = (~t[255] & t[256]);
  assign t[20] = t[30] ^ t[31];
  assign t[210] = (~t[257] & t[258]);
  assign t[211] = (~t[259] & t[260]);
  assign t[212] = (~t[261] & t[262]);
  assign t[213] = (~t[263] & t[264]);
  assign t[214] = (~t[265] & t[266]);
  assign t[215] = (~t[263] & t[267]);
  assign t[216] = (~t[263] & t[268]);
  assign t[217] = (~t[269] & t[270]);
  assign t[218] = (~t[271] & t[272]);
  assign t[219] = (~t[273] & t[274]);
  assign t[21] = x[7] ? t[33] : t[32];
  assign t[220] = (~t[265] & t[275]);
  assign t[221] = (~t[265] & t[276]);
  assign t[222] = (~t[277] & t[278]);
  assign t[223] = (~t[279] & t[280]);
  assign t[224] = (~t[281] & t[282]);
  assign t[225] = (~t[263] & t[283]);
  assign t[226] = (~t[269] & t[284]);
  assign t[227] = (~t[269] & t[285]);
  assign t[228] = (~t[271] & t[286]);
  assign t[229] = (~t[271] & t[287]);
  assign t[22] = x[7] ? t[35] : t[34];
  assign t[230] = (~t[273] & t[288]);
  assign t[231] = (~t[273] & t[289]);
  assign t[232] = (~t[265] & t[290]);
  assign t[233] = (~t[277] & t[291]);
  assign t[234] = (~t[277] & t[292]);
  assign t[235] = (~t[279] & t[293]);
  assign t[236] = (~t[279] & t[294]);
  assign t[237] = (~t[295] & t[296]);
  assign t[238] = (~t[281] & t[297]);
  assign t[239] = (~t[281] & t[298]);
  assign t[23] = ~(t[121]);
  assign t[240] = (~t[299] & t[300]);
  assign t[241] = (~t[269] & t[301]);
  assign t[242] = (~t[271] & t[302]);
  assign t[243] = (~t[273] & t[303]);
  assign t[244] = (~t[277] & t[304]);
  assign t[245] = (~t[279] & t[305]);
  assign t[246] = (~t[295] & t[306]);
  assign t[247] = (~t[295] & t[307]);
  assign t[248] = (~t[281] & t[308]);
  assign t[249] = (~t[299] & t[309]);
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = (~t[299] & t[310]);
  assign t[251] = (~t[295] & t[311]);
  assign t[252] = (~t[299] & t[312]);
  assign t[253] = t[313] ^ x[4];
  assign t[254] = t[314] ^ x[5];
  assign t[255] = t[315] ^ x[10];
  assign t[256] = t[316] ^ x[11];
  assign t[257] = t[317] ^ x[13];
  assign t[258] = t[318] ^ x[14];
  assign t[259] = t[319] ^ x[16];
  assign t[25] = t[38] ^ t[39];
  assign t[260] = t[320] ^ x[17];
  assign t[261] = t[321] ^ x[19];
  assign t[262] = t[322] ^ x[20];
  assign t[263] = t[323] ^ x[27];
  assign t[264] = t[324] ^ x[28];
  assign t[265] = t[325] ^ x[35];
  assign t[266] = t[326] ^ x[36];
  assign t[267] = t[327] ^ x[39];
  assign t[268] = t[328] ^ x[40];
  assign t[269] = t[329] ^ x[45];
  assign t[26] = x[7] ? t[41] : t[40];
  assign t[270] = t[330] ^ x[46];
  assign t[271] = t[331] ^ x[51];
  assign t[272] = t[332] ^ x[52];
  assign t[273] = t[333] ^ x[59];
  assign t[274] = t[334] ^ x[60];
  assign t[275] = t[335] ^ x[63];
  assign t[276] = t[336] ^ x[64];
  assign t[277] = t[337] ^ x[69];
  assign t[278] = t[338] ^ x[70];
  assign t[279] = t[339] ^ x[75];
  assign t[27] = x[7] ? t[43] : t[42];
  assign t[280] = t[340] ^ x[76];
  assign t[281] = t[341] ^ x[83];
  assign t[282] = t[342] ^ x[84];
  assign t[283] = t[343] ^ x[87];
  assign t[284] = t[344] ^ x[88];
  assign t[285] = t[345] ^ x[89];
  assign t[286] = t[346] ^ x[90];
  assign t[287] = t[347] ^ x[91];
  assign t[288] = t[348] ^ x[92];
  assign t[289] = t[349] ^ x[93];
  assign t[28] = ~(t[44] & t[45]);
  assign t[290] = t[350] ^ x[94];
  assign t[291] = t[351] ^ x[95];
  assign t[292] = t[352] ^ x[96];
  assign t[293] = t[353] ^ x[97];
  assign t[294] = t[354] ^ x[98];
  assign t[295] = t[355] ^ x[103];
  assign t[296] = t[356] ^ x[104];
  assign t[297] = t[357] ^ x[105];
  assign t[298] = t[358] ^ x[106];
  assign t[299] = t[359] ^ x[111];
  assign t[29] = ~(t[46] & t[123]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = t[360] ^ x[112];
  assign t[301] = t[361] ^ x[113];
  assign t[302] = t[362] ^ x[114];
  assign t[303] = t[363] ^ x[115];
  assign t[304] = t[364] ^ x[116];
  assign t[305] = t[365] ^ x[117];
  assign t[306] = t[366] ^ x[118];
  assign t[307] = t[367] ^ x[119];
  assign t[308] = t[368] ^ x[120];
  assign t[309] = t[369] ^ x[121];
  assign t[30] = t[16] ? x[30] : x[29];
  assign t[310] = t[370] ^ x[122];
  assign t[311] = t[371] ^ x[123];
  assign t[312] = t[372] ^ x[124];
  assign t[313] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[314] = (x[2]);
  assign t[315] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[316] = (x[9]);
  assign t[317] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[318] = (x[12]);
  assign t[319] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = ~(t[47] & t[48]);
  assign t[320] = (x[15]);
  assign t[321] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[322] = (x[18]);
  assign t[323] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[324] = (x[24]);
  assign t[325] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[326] = (x[32]);
  assign t[327] = (x[26]);
  assign t[328] = (x[23]);
  assign t[329] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[32] = ~(t[49] & t[50]);
  assign t[330] = (x[42]);
  assign t[331] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[332] = (x[48]);
  assign t[333] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[334] = (x[56]);
  assign t[335] = (x[34]);
  assign t[336] = (x[31]);
  assign t[337] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[338] = (x[66]);
  assign t[339] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[33] = t[51] ^ t[32];
  assign t[340] = (x[72]);
  assign t[341] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[342] = (x[80]);
  assign t[343] = (x[25]);
  assign t[344] = (x[44]);
  assign t[345] = (x[41]);
  assign t[346] = (x[50]);
  assign t[347] = (x[47]);
  assign t[348] = (x[58]);
  assign t[349] = (x[55]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[33]);
  assign t[351] = (x[68]);
  assign t[352] = (x[65]);
  assign t[353] = (x[74]);
  assign t[354] = (x[71]);
  assign t[355] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[356] = (x[100]);
  assign t[357] = (x[82]);
  assign t[358] = (x[79]);
  assign t[359] = (x[107] & ~x[108] & ~x[109] & ~x[110]) | (~x[107] & x[108] & ~x[109] & ~x[110]) | (~x[107] & ~x[108] & x[109] & ~x[110]) | (~x[107] & ~x[108] & ~x[109] & x[110]) | (x[107] & x[108] & x[109] & ~x[110]) | (x[107] & x[108] & ~x[109] & x[110]) | (x[107] & ~x[108] & x[109] & x[110]) | (~x[107] & x[108] & x[109] & x[110]);
  assign t[35] = t[54] ^ t[40];
  assign t[360] = (x[108]);
  assign t[361] = (x[43]);
  assign t[362] = (x[49]);
  assign t[363] = (x[57]);
  assign t[364] = (x[67]);
  assign t[365] = (x[73]);
  assign t[366] = (x[102]);
  assign t[367] = (x[99]);
  assign t[368] = (x[81]);
  assign t[369] = (x[110]);
  assign t[36] = ~(t[55] & t[56]);
  assign t[370] = (x[107]);
  assign t[371] = (x[101]);
  assign t[372] = (x[109]);
  assign t[37] = ~(t[57] & t[124]);
  assign t[38] = t[16] ? x[38] : x[37];
  assign t[39] = ~(t[58] & t[59]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[60] & t[61]);
  assign t[41] = t[62] ^ t[63];
  assign t[42] = ~(t[64] & t[65]);
  assign t[43] = t[66] ^ t[67];
  assign t[44] = ~(t[125]);
  assign t[45] = ~(t[126]);
  assign t[46] = ~(t[68] & t[69]);
  assign t[47] = ~(t[70] & t[71]);
  assign t[48] = ~(t[72] & t[127]);
  assign t[49] = ~(t[73] & t[74]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[75] & t[128]);
  assign t[51] = t[76] ? x[54] : x[53];
  assign t[52] = ~(t[77] & t[78]);
  assign t[53] = ~(t[79] & t[129]);
  assign t[54] = t[76] ? x[62] : x[61];
  assign t[55] = ~(t[130]);
  assign t[56] = ~(t[131]);
  assign t[57] = ~(t[80] & t[81]);
  assign t[58] = ~(t[82] & t[83]);
  assign t[59] = ~(t[84] & t[132]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[85] & t[86]);
  assign t[61] = ~(t[87] & t[133]);
  assign t[62] = t[88] ? x[78] : x[77];
  assign t[63] = ~(t[89] & t[90]);
  assign t[64] = ~(t[91] & t[92]);
  assign t[65] = ~(t[93] & t[134]);
  assign t[66] = t[88] ? x[86] : x[85];
  assign t[67] = ~(t[94] & t[95]);
  assign t[68] = ~(t[126] & t[125]);
  assign t[69] = ~(t[135]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[136]);
  assign t[71] = ~(t[137]);
  assign t[72] = ~(t[96] & t[97]);
  assign t[73] = ~(t[138]);
  assign t[74] = ~(t[139]);
  assign t[75] = ~(t[98] & t[99]);
  assign t[76] = ~(t[23]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = ~(t[119] & t[120]);
  assign t[80] = ~(t[131] & t[130]);
  assign t[81] = ~(t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[102] & t[103]);
  assign t[85] = ~(t[145]);
  assign t[86] = ~(t[146]);
  assign t[87] = ~(t[104] & t[105]);
  assign t[88] = ~(t[23]);
  assign t[89] = ~(t[106] & t[107]);
  assign t[8] = ~(t[121] & t[122]);
  assign t[90] = ~(t[108] & t[147]);
  assign t[91] = ~(t[148]);
  assign t[92] = ~(t[149]);
  assign t[93] = ~(t[109] & t[110]);
  assign t[94] = ~(t[111] & t[112]);
  assign t[95] = ~(t[113] & t[150]);
  assign t[96] = ~(t[137] & t[136]);
  assign t[97] = ~(t[151]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[152]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [114:0] x;
 output y;

 wire [302:0] t;
  assign t[0] = t[1] ? t[2] : t[98];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[14] ^ t[15]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = x[21] ^ x[22];
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[16] ? x[22] : x[21];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = t[168] ^ x[5];
  assign t[134] = t[169] ^ x[11];
  assign t[135] = t[170] ^ x[14];
  assign t[136] = t[171] ^ x[17];
  assign t[137] = t[172] ^ x[20];
  assign t[138] = t[173] ^ x[28];
  assign t[139] = t[174] ^ x[29];
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = t[175] ^ x[37];
  assign t[141] = t[176] ^ x[38];
  assign t[142] = t[177] ^ x[41];
  assign t[143] = t[178] ^ x[47];
  assign t[144] = t[179] ^ x[48];
  assign t[145] = t[180] ^ x[54];
  assign t[146] = t[181] ^ x[55];
  assign t[147] = t[182] ^ x[63];
  assign t[148] = t[183] ^ x[64];
  assign t[149] = t[184] ^ x[67];
  assign t[14] = x[7] ? t[20] : t[19];
  assign t[150] = t[185] ^ x[73];
  assign t[151] = t[186] ^ x[74];
  assign t[152] = t[187] ^ x[80];
  assign t[153] = t[188] ^ x[81];
  assign t[154] = t[189] ^ x[89];
  assign t[155] = t[190] ^ x[90];
  assign t[156] = t[191] ^ x[93];
  assign t[157] = t[192] ^ x[94];
  assign t[158] = t[193] ^ x[95];
  assign t[159] = t[194] ^ x[96];
  assign t[15] = ~(t[21] ^ t[22]);
  assign t[160] = t[195] ^ x[97];
  assign t[161] = t[196] ^ x[103];
  assign t[162] = t[197] ^ x[104];
  assign t[163] = t[198] ^ x[105];
  assign t[164] = t[199] ^ x[111];
  assign t[165] = t[200] ^ x[112];
  assign t[166] = t[201] ^ x[113];
  assign t[167] = t[202] ^ x[114];
  assign t[168] = (~t[203] & t[204]);
  assign t[169] = (~t[205] & t[206]);
  assign t[16] = ~(t[23]);
  assign t[170] = (~t[207] & t[208]);
  assign t[171] = (~t[209] & t[210]);
  assign t[172] = (~t[211] & t[212]);
  assign t[173] = (~t[213] & t[214]);
  assign t[174] = (~t[213] & t[215]);
  assign t[175] = (~t[216] & t[217]);
  assign t[176] = (~t[216] & t[218]);
  assign t[177] = (~t[213] & t[219]);
  assign t[178] = (~t[220] & t[221]);
  assign t[179] = (~t[220] & t[222]);
  assign t[17] = x[7] ? t[25] : t[24];
  assign t[180] = (~t[223] & t[224]);
  assign t[181] = (~t[223] & t[225]);
  assign t[182] = (~t[226] & t[227]);
  assign t[183] = (~t[226] & t[228]);
  assign t[184] = (~t[216] & t[229]);
  assign t[185] = (~t[230] & t[231]);
  assign t[186] = (~t[230] & t[232]);
  assign t[187] = (~t[233] & t[234]);
  assign t[188] = (~t[233] & t[235]);
  assign t[189] = (~t[236] & t[237]);
  assign t[18] = ~(t[26] ^ t[27]);
  assign t[190] = (~t[236] & t[238]);
  assign t[191] = (~t[220] & t[239]);
  assign t[192] = (~t[223] & t[240]);
  assign t[193] = (~t[226] & t[241]);
  assign t[194] = (~t[230] & t[242]);
  assign t[195] = (~t[233] & t[243]);
  assign t[196] = (~t[244] & t[245]);
  assign t[197] = (~t[244] & t[246]);
  assign t[198] = (~t[236] & t[247]);
  assign t[199] = (~t[248] & t[249]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = (~t[248] & t[250]);
  assign t[201] = (~t[244] & t[251]);
  assign t[202] = (~t[248] & t[252]);
  assign t[203] = t[253] ^ x[4];
  assign t[204] = t[254] ^ x[5];
  assign t[205] = t[255] ^ x[10];
  assign t[206] = t[256] ^ x[11];
  assign t[207] = t[257] ^ x[13];
  assign t[208] = t[258] ^ x[14];
  assign t[209] = t[259] ^ x[16];
  assign t[20] = t[30] ^ t[31];
  assign t[210] = t[260] ^ x[17];
  assign t[211] = t[261] ^ x[19];
  assign t[212] = t[262] ^ x[20];
  assign t[213] = t[263] ^ x[27];
  assign t[214] = t[264] ^ x[28];
  assign t[215] = t[265] ^ x[29];
  assign t[216] = t[266] ^ x[36];
  assign t[217] = t[267] ^ x[37];
  assign t[218] = t[268] ^ x[38];
  assign t[219] = t[269] ^ x[41];
  assign t[21] = x[7] ? t[33] : t[32];
  assign t[220] = t[270] ^ x[46];
  assign t[221] = t[271] ^ x[47];
  assign t[222] = t[272] ^ x[48];
  assign t[223] = t[273] ^ x[53];
  assign t[224] = t[274] ^ x[54];
  assign t[225] = t[275] ^ x[55];
  assign t[226] = t[276] ^ x[62];
  assign t[227] = t[277] ^ x[63];
  assign t[228] = t[278] ^ x[64];
  assign t[229] = t[279] ^ x[67];
  assign t[22] = x[7] ? t[35] : t[34];
  assign t[230] = t[280] ^ x[72];
  assign t[231] = t[281] ^ x[73];
  assign t[232] = t[282] ^ x[74];
  assign t[233] = t[283] ^ x[79];
  assign t[234] = t[284] ^ x[80];
  assign t[235] = t[285] ^ x[81];
  assign t[236] = t[286] ^ x[88];
  assign t[237] = t[287] ^ x[89];
  assign t[238] = t[288] ^ x[90];
  assign t[239] = t[289] ^ x[93];
  assign t[23] = ~(t[101]);
  assign t[240] = t[290] ^ x[94];
  assign t[241] = t[291] ^ x[95];
  assign t[242] = t[292] ^ x[96];
  assign t[243] = t[293] ^ x[97];
  assign t[244] = t[294] ^ x[102];
  assign t[245] = t[295] ^ x[103];
  assign t[246] = t[296] ^ x[104];
  assign t[247] = t[297] ^ x[105];
  assign t[248] = t[298] ^ x[110];
  assign t[249] = t[299] ^ x[111];
  assign t[24] = ~(t[36] & t[37]);
  assign t[250] = t[300] ^ x[112];
  assign t[251] = t[301] ^ x[113];
  assign t[252] = t[302] ^ x[114];
  assign t[253] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[254] = (x[1]);
  assign t[255] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[256] = (x[9]);
  assign t[257] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[258] = (x[12]);
  assign t[259] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[25] = t[38] ^ t[39];
  assign t[260] = (x[15]);
  assign t[261] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[262] = (x[18]);
  assign t[263] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[264] = (x[25]);
  assign t[265] = (x[23]);
  assign t[266] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[267] = (x[34]);
  assign t[268] = (x[32]);
  assign t[269] = (x[26]);
  assign t[26] = x[7] ? t[41] : t[40];
  assign t[270] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[271] = (x[44]);
  assign t[272] = (x[42]);
  assign t[273] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[274] = (x[51]);
  assign t[275] = (x[49]);
  assign t[276] = (x[58] & ~x[59] & ~x[60] & ~x[61]) | (~x[58] & x[59] & ~x[60] & ~x[61]) | (~x[58] & ~x[59] & x[60] & ~x[61]) | (~x[58] & ~x[59] & ~x[60] & x[61]) | (x[58] & x[59] & x[60] & ~x[61]) | (x[58] & x[59] & ~x[60] & x[61]) | (x[58] & ~x[59] & x[60] & x[61]) | (~x[58] & x[59] & x[60] & x[61]);
  assign t[277] = (x[60]);
  assign t[278] = (x[58]);
  assign t[279] = (x[35]);
  assign t[27] = x[7] ? t[43] : t[42];
  assign t[280] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[281] = (x[70]);
  assign t[282] = (x[68]);
  assign t[283] = (x[75] & ~x[76] & ~x[77] & ~x[78]) | (~x[75] & x[76] & ~x[77] & ~x[78]) | (~x[75] & ~x[76] & x[77] & ~x[78]) | (~x[75] & ~x[76] & ~x[77] & x[78]) | (x[75] & x[76] & x[77] & ~x[78]) | (x[75] & x[76] & ~x[77] & x[78]) | (x[75] & ~x[76] & x[77] & x[78]) | (~x[75] & x[76] & x[77] & x[78]);
  assign t[284] = (x[77]);
  assign t[285] = (x[75]);
  assign t[286] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[287] = (x[86]);
  assign t[288] = (x[84]);
  assign t[289] = (x[45]);
  assign t[28] = ~(t[103] & t[44]);
  assign t[290] = (x[52]);
  assign t[291] = (x[61]);
  assign t[292] = (x[71]);
  assign t[293] = (x[78]);
  assign t[294] = (x[98] & ~x[99] & ~x[100] & ~x[101]) | (~x[98] & x[99] & ~x[100] & ~x[101]) | (~x[98] & ~x[99] & x[100] & ~x[101]) | (~x[98] & ~x[99] & ~x[100] & x[101]) | (x[98] & x[99] & x[100] & ~x[101]) | (x[98] & x[99] & ~x[100] & x[101]) | (x[98] & ~x[99] & x[100] & x[101]) | (~x[98] & x[99] & x[100] & x[101]);
  assign t[295] = (x[100]);
  assign t[296] = (x[98]);
  assign t[297] = (x[87]);
  assign t[298] = (x[106] & ~x[107] & ~x[108] & ~x[109]) | (~x[106] & x[107] & ~x[108] & ~x[109]) | (~x[106] & ~x[107] & x[108] & ~x[109]) | (~x[106] & ~x[107] & ~x[108] & x[109]) | (x[106] & x[107] & x[108] & ~x[109]) | (x[106] & x[107] & ~x[108] & x[109]) | (x[106] & ~x[107] & x[108] & x[109]) | (~x[106] & x[107] & x[108] & x[109]);
  assign t[299] = (x[108]);
  assign t[29] = ~(t[104] & t[45]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[300] = (x[106]);
  assign t[301] = (x[101]);
  assign t[302] = (x[109]);
  assign t[30] = t[16] ? x[31] : x[30];
  assign t[31] = ~(t[46] & t[47]);
  assign t[32] = ~(t[48] & t[49]);
  assign t[33] = t[50] ^ t[40];
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[34];
  assign t[36] = ~(t[105] & t[54]);
  assign t[37] = ~(t[106] & t[55]);
  assign t[38] = t[16] ? x[40] : x[39];
  assign t[39] = ~(t[56] & t[57]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[58] & t[59]);
  assign t[41] = t[60] ^ t[61];
  assign t[42] = ~(t[62] & t[63]);
  assign t[43] = t[64] ^ t[65];
  assign t[44] = ~(t[107]);
  assign t[45] = ~(t[107] & t[66]);
  assign t[46] = ~(t[108] & t[67]);
  assign t[47] = ~(t[109] & t[68]);
  assign t[48] = ~(t[110] & t[69]);
  assign t[49] = ~(t[111] & t[70]);
  assign t[4] = ~(x[6]);
  assign t[50] = t[71] ? x[57] : x[56];
  assign t[51] = ~(t[112] & t[72]);
  assign t[52] = ~(t[113] & t[73]);
  assign t[53] = t[71] ? x[66] : x[65];
  assign t[54] = ~(t[114]);
  assign t[55] = ~(t[114] & t[74]);
  assign t[56] = ~(t[115] & t[75]);
  assign t[57] = ~(t[116] & t[76]);
  assign t[58] = ~(t[117] & t[77]);
  assign t[59] = ~(t[118] & t[78]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[79] ? x[83] : x[82];
  assign t[61] = ~(t[80] & t[81]);
  assign t[62] = ~(t[119] & t[82]);
  assign t[63] = ~(t[120] & t[83]);
  assign t[64] = t[79] ? x[92] : x[91];
  assign t[65] = ~(t[84] & t[85]);
  assign t[66] = ~(t[103]);
  assign t[67] = ~(t[121]);
  assign t[68] = ~(t[121] & t[86]);
  assign t[69] = ~(t[122]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[122] & t[87]);
  assign t[71] = ~(t[23]);
  assign t[72] = ~(t[123]);
  assign t[73] = ~(t[123] & t[88]);
  assign t[74] = ~(t[105]);
  assign t[75] = ~(t[124]);
  assign t[76] = ~(t[124] & t[89]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[125] & t[90]);
  assign t[79] = ~(t[23]);
  assign t[7] = ~(t[99] & t[100]);
  assign t[80] = ~(t[126] & t[91]);
  assign t[81] = ~(t[127] & t[92]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[128] & t[93]);
  assign t[84] = ~(t[129] & t[94]);
  assign t[85] = ~(t[130] & t[95]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[112]);
  assign t[89] = ~(t[115]);
  assign t[8] = ~(t[101] & t[102]);
  assign t[90] = ~(t[117]);
  assign t[91] = ~(t[131]);
  assign t[92] = ~(t[131] & t[96]);
  assign t[93] = ~(t[119]);
  assign t[94] = ~(t[132]);
  assign t[95] = ~(t[132] & t[97]);
  assign t[96] = ~(t[126]);
  assign t[97] = ~(t[129]);
  assign t[98] = (t[133]);
  assign t[99] = (t[134]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [124:0] x;
 output y;

 wire [455:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = t[135] ? x[89] : x[88];
  assign t[101] = ~(t[139] & t[140]);
  assign t[102] = ~(t[225]);
  assign t[103] = ~(t[213] | t[214]);
  assign t[104] = ~(t[226]);
  assign t[105] = ~(t[227]);
  assign t[106] = ~(t[141] | t[142]);
  assign t[107] = ~(t[139] & t[143]);
  assign t[108] = ~(t[228]);
  assign t[109] = ~(t[229]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[144] | t[145]);
  assign t[111] = ~(t[146] | t[147]);
  assign t[112] = ~(t[230] | t[148]);
  assign t[113] = t[149] ? x[102] : x[101];
  assign t[114] = ~(t[150] & t[151]);
  assign t[115] = ~(t[231]);
  assign t[116] = ~(t[232]);
  assign t[117] = ~(t[152] | t[153]);
  assign t[118] = ~(t[154] | t[155]);
  assign t[119] = ~(t[233] | t[156]);
  assign t[11] = ~(x[6]);
  assign t[120] = t[149] ? x[112] : x[111];
  assign t[121] = ~(t[157] & t[143]);
  assign t[122] = ~(t[204]);
  assign t[123] = ~(t[158] & t[159]);
  assign t[124] = ~(t[160] & t[205]);
  assign t[125] = ~(t[81] | t[161]);
  assign t[126] = ~(t[81] | t[162]);
  assign t[127] = ~(x[7] & t[163]);
  assign t[128] = ~(t[205] & t[164]);
  assign t[129] = ~(t[234]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[219] | t[220]);
  assign t[131] = ~(t[157] & t[139]);
  assign t[132] = ~(t[81] | t[165]);
  assign t[133] = ~(t[235]);
  assign t[134] = ~(t[221] | t[222]);
  assign t[135] = ~(t[49]);
  assign t[136] = ~(t[166] | t[167]);
  assign t[137] = ~(t[236]);
  assign t[138] = ~(t[223] | t[224]);
  assign t[139] = ~(t[168] | t[167]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[169] | t[170]);
  assign t[141] = ~(t[237]);
  assign t[142] = ~(t[226] | t[227]);
  assign t[143] = ~(t[171] & t[172]);
  assign t[144] = ~(t[238]);
  assign t[145] = ~(t[228] | t[229]);
  assign t[146] = ~(t[239]);
  assign t[147] = ~(t[240]);
  assign t[148] = ~(t[173] | t[174]);
  assign t[149] = ~(t[49]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[175] | t[176]);
  assign t[151] = ~(t[177] & t[178]);
  assign t[152] = ~(t[241]);
  assign t[153] = ~(t[231] | t[232]);
  assign t[154] = ~(t[242]);
  assign t[155] = ~(t[243]);
  assign t[156] = ~(t[179] | t[180]);
  assign t[157] = ~(t[50] | t[169]);
  assign t[158] = ~(x[7] | t[203]);
  assign t[159] = ~(t[205]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = x[7] & t[203];
  assign t[161] = t[202] ? t[182] : t[181];
  assign t[162] = t[202] ? t[184] : t[183];
  assign t[163] = ~(t[203] | t[205]);
  assign t[164] = ~(x[7] | t[185]);
  assign t[165] = t[202] ? t[123] : t[124];
  assign t[166] = ~(t[122] | t[186]);
  assign t[167] = ~(t[122] | t[187]);
  assign t[168] = ~(t[122] | t[188]);
  assign t[169] = ~(t[189] & t[190]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[151] & t[191]);
  assign t[171] = ~(t[203] | t[159]);
  assign t[172] = t[81] & t[202];
  assign t[173] = ~(t[244]);
  assign t[174] = ~(t[239] | t[240]);
  assign t[175] = ~(t[192] & t[143]);
  assign t[176] = t[52] | t[193];
  assign t[177] = t[205] & t[194];
  assign t[178] = t[158] | t[160];
  assign t[179] = ~(t[245]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[242] | t[243]);
  assign t[181] = ~(t[164] & t[159]);
  assign t[182] = ~(x[7] & t[171]);
  assign t[183] = ~(t[158] & t[205]);
  assign t[184] = ~(t[160] & t[159]);
  assign t[185] = ~(t[203]);
  assign t[186] = t[202] ? t[123] : t[184];
  assign t[187] = t[202] ? t[181] : t[127];
  assign t[188] = t[202] ? t[184] : t[123];
  assign t[189] = ~(t[166] | t[195]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[122] & t[196]);
  assign t[191] = t[122] | t[197];
  assign t[192] = ~(t[194] & t[198]);
  assign t[193] = ~(t[81] | t[199]);
  assign t[194] = ~(t[122] | t[202]);
  assign t[195] = ~(t[81] | t[200]);
  assign t[196] = ~(t[127] & t[128]);
  assign t[197] = t[202] ? t[127] : t[181];
  assign t[198] = ~(t[128] & t[182]);
  assign t[199] = t[202] ? t[183] : t[184];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[181] : t[182];
  assign t[201] = (t[246]);
  assign t[202] = (t[247]);
  assign t[203] = (t[248]);
  assign t[204] = (t[249]);
  assign t[205] = (t[250]);
  assign t[206] = (t[251]);
  assign t[207] = (t[252]);
  assign t[208] = (t[253]);
  assign t[209] = (t[254]);
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = (t[255]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = t[291] ^ x[5];
  assign t[247] = t[292] ^ x[13];
  assign t[248] = t[293] ^ x[16];
  assign t[249] = t[294] ^ x[19];
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = t[295] ^ x[22];
  assign t[251] = t[296] ^ x[28];
  assign t[252] = t[297] ^ x[34];
  assign t[253] = t[298] ^ x[35];
  assign t[254] = t[299] ^ x[36];
  assign t[255] = t[300] ^ x[42];
  assign t[256] = t[301] ^ x[50];
  assign t[257] = t[302] ^ x[56];
  assign t[258] = t[303] ^ x[57];
  assign t[259] = t[304] ^ x[58];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[64];
  assign t[261] = t[306] ^ x[72];
  assign t[262] = t[307] ^ x[78];
  assign t[263] = t[308] ^ x[79];
  assign t[264] = t[309] ^ x[80];
  assign t[265] = t[310] ^ x[81];
  assign t[266] = t[311] ^ x[82];
  assign t[267] = t[312] ^ x[83];
  assign t[268] = t[313] ^ x[86];
  assign t[269] = t[314] ^ x[87];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[90];
  assign t[271] = t[316] ^ x[91];
  assign t[272] = t[317] ^ x[92];
  assign t[273] = t[318] ^ x[93];
  assign t[274] = t[319] ^ x[94];
  assign t[275] = t[320] ^ x[100];
  assign t[276] = t[321] ^ x[103];
  assign t[277] = t[322] ^ x[104];
  assign t[278] = t[323] ^ x[110];
  assign t[279] = t[324] ^ x[113];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[114];
  assign t[281] = t[326] ^ x[115];
  assign t[282] = t[327] ^ x[116];
  assign t[283] = t[328] ^ x[117];
  assign t[284] = t[329] ^ x[118];
  assign t[285] = t[330] ^ x[119];
  assign t[286] = t[331] ^ x[120];
  assign t[287] = t[332] ^ x[121];
  assign t[288] = t[333] ^ x[122];
  assign t[289] = t[334] ^ x[123];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[124];
  assign t[291] = (~t[336] & t[337]);
  assign t[292] = (~t[338] & t[339]);
  assign t[293] = (~t[340] & t[341]);
  assign t[294] = (~t[342] & t[343]);
  assign t[295] = (~t[344] & t[345]);
  assign t[296] = (~t[346] & t[347]);
  assign t[297] = (~t[348] & t[349]);
  assign t[298] = (~t[346] & t[350]);
  assign t[299] = (~t[346] & t[351]);
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[352] & t[353]);
  assign t[301] = (~t[354] & t[355]);
  assign t[302] = (~t[356] & t[357]);
  assign t[303] = (~t[348] & t[358]);
  assign t[304] = (~t[348] & t[359]);
  assign t[305] = (~t[360] & t[361]);
  assign t[306] = (~t[362] & t[363]);
  assign t[307] = (~t[364] & t[365]);
  assign t[308] = (~t[346] & t[366]);
  assign t[309] = (~t[352] & t[367]);
  assign t[30] = ~(t[49]);
  assign t[310] = (~t[352] & t[368]);
  assign t[311] = (~t[354] & t[369]);
  assign t[312] = (~t[354] & t[370]);
  assign t[313] = (~t[356] & t[371]);
  assign t[314] = (~t[356] & t[372]);
  assign t[315] = (~t[348] & t[373]);
  assign t[316] = (~t[360] & t[374]);
  assign t[317] = (~t[360] & t[375]);
  assign t[318] = (~t[362] & t[376]);
  assign t[319] = (~t[362] & t[377]);
  assign t[31] = ~(t[50]);
  assign t[320] = (~t[378] & t[379]);
  assign t[321] = (~t[364] & t[380]);
  assign t[322] = (~t[364] & t[381]);
  assign t[323] = (~t[382] & t[383]);
  assign t[324] = (~t[352] & t[384]);
  assign t[325] = (~t[354] & t[385]);
  assign t[326] = (~t[356] & t[386]);
  assign t[327] = (~t[360] & t[387]);
  assign t[328] = (~t[362] & t[388]);
  assign t[329] = (~t[378] & t[389]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = (~t[378] & t[390]);
  assign t[331] = (~t[364] & t[391]);
  assign t[332] = (~t[382] & t[392]);
  assign t[333] = (~t[382] & t[393]);
  assign t[334] = (~t[378] & t[394]);
  assign t[335] = (~t[382] & t[395]);
  assign t[336] = t[396] ^ x[4];
  assign t[337] = t[397] ^ x[5];
  assign t[338] = t[398] ^ x[12];
  assign t[339] = t[399] ^ x[13];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[400] ^ x[15];
  assign t[341] = t[401] ^ x[16];
  assign t[342] = t[402] ^ x[18];
  assign t[343] = t[403] ^ x[19];
  assign t[344] = t[404] ^ x[21];
  assign t[345] = t[405] ^ x[22];
  assign t[346] = t[406] ^ x[27];
  assign t[347] = t[407] ^ x[28];
  assign t[348] = t[408] ^ x[33];
  assign t[349] = t[409] ^ x[34];
  assign t[34] = ~(t[206] | t[55]);
  assign t[350] = t[410] ^ x[35];
  assign t[351] = t[411] ^ x[36];
  assign t[352] = t[412] ^ x[41];
  assign t[353] = t[413] ^ x[42];
  assign t[354] = t[414] ^ x[49];
  assign t[355] = t[415] ^ x[50];
  assign t[356] = t[416] ^ x[55];
  assign t[357] = t[417] ^ x[56];
  assign t[358] = t[418] ^ x[57];
  assign t[359] = t[419] ^ x[58];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[420] ^ x[63];
  assign t[361] = t[421] ^ x[64];
  assign t[362] = t[422] ^ x[71];
  assign t[363] = t[423] ^ x[72];
  assign t[364] = t[424] ^ x[77];
  assign t[365] = t[425] ^ x[78];
  assign t[366] = t[426] ^ x[79];
  assign t[367] = t[427] ^ x[80];
  assign t[368] = t[428] ^ x[81];
  assign t[369] = t[429] ^ x[82];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[430] ^ x[83];
  assign t[371] = t[431] ^ x[86];
  assign t[372] = t[432] ^ x[87];
  assign t[373] = t[433] ^ x[90];
  assign t[374] = t[434] ^ x[91];
  assign t[375] = t[435] ^ x[92];
  assign t[376] = t[436] ^ x[93];
  assign t[377] = t[437] ^ x[94];
  assign t[378] = t[438] ^ x[99];
  assign t[379] = t[439] ^ x[100];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[440] ^ x[103];
  assign t[381] = t[441] ^ x[104];
  assign t[382] = t[442] ^ x[109];
  assign t[383] = t[443] ^ x[110];
  assign t[384] = t[444] ^ x[113];
  assign t[385] = t[445] ^ x[114];
  assign t[386] = t[446] ^ x[115];
  assign t[387] = t[447] ^ x[116];
  assign t[388] = t[448] ^ x[117];
  assign t[389] = t[449] ^ x[118];
  assign t[38] = ~(t[37] ^ t[62]);
  assign t[390] = t[450] ^ x[119];
  assign t[391] = t[451] ^ x[120];
  assign t[392] = t[452] ^ x[121];
  assign t[393] = t[453] ^ x[122];
  assign t[394] = t[454] ^ x[123];
  assign t[395] = t[455] ^ x[124];
  assign t[396] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[397] = (x[0]);
  assign t[398] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[399] = (x[11]);
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[401] = (x[14]);
  assign t[402] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[403] = (x[17]);
  assign t[404] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[405] = (x[20]);
  assign t[406] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[407] = (x[24]);
  assign t[408] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[409] = (x[30]);
  assign t[40] = ~(t[47] ^ t[65]);
  assign t[410] = (x[25]);
  assign t[411] = (x[26]);
  assign t[412] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[413] = (x[38]);
  assign t[414] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[415] = (x[46]);
  assign t[416] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[417] = (x[52]);
  assign t[418] = (x[31]);
  assign t[419] = (x[32]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[421] = (x[60]);
  assign t[422] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[423] = (x[68]);
  assign t[424] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[425] = (x[74]);
  assign t[426] = (x[23]);
  assign t[427] = (x[39]);
  assign t[428] = (x[40]);
  assign t[429] = (x[47]);
  assign t[42] = ~(t[207] | t[68]);
  assign t[430] = (x[48]);
  assign t[431] = (x[53]);
  assign t[432] = (x[54]);
  assign t[433] = (x[29]);
  assign t[434] = (x[61]);
  assign t[435] = (x[62]);
  assign t[436] = (x[69]);
  assign t[437] = (x[70]);
  assign t[438] = (x[95] & ~x[96] & ~x[97] & ~x[98]) | (~x[95] & x[96] & ~x[97] & ~x[98]) | (~x[95] & ~x[96] & x[97] & ~x[98]) | (~x[95] & ~x[96] & ~x[97] & x[98]) | (x[95] & x[96] & x[97] & ~x[98]) | (x[95] & x[96] & ~x[97] & x[98]) | (x[95] & ~x[96] & x[97] & x[98]) | (~x[95] & x[96] & x[97] & x[98]);
  assign t[439] = (x[96]);
  assign t[43] = ~(t[69] | t[70]);
  assign t[440] = (x[75]);
  assign t[441] = (x[76]);
  assign t[442] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[443] = (x[106]);
  assign t[444] = (x[37]);
  assign t[445] = (x[45]);
  assign t[446] = (x[51]);
  assign t[447] = (x[59]);
  assign t[448] = (x[67]);
  assign t[449] = (x[97]);
  assign t[44] = ~(t[71] ^ t[72]);
  assign t[450] = (x[98]);
  assign t[451] = (x[73]);
  assign t[452] = (x[107]);
  assign t[453] = (x[108]);
  assign t[454] = (x[95]);
  assign t[455] = (x[105]);
  assign t[45] = ~(t[73] | t[74]);
  assign t[46] = ~(t[75] ^ t[76]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[48] = ~(t[79] ^ t[80]);
  assign t[49] = ~(t[204]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[81] | t[82]);
  assign t[51] = ~(t[83]);
  assign t[52] = ~(t[81] | t[84]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[209]);
  assign t[55] = ~(t[85] | t[86]);
  assign t[56] = ~(t[87] | t[88]);
  assign t[57] = ~(t[210] | t[89]);
  assign t[58] = t[30] ? x[44] : x[43];
  assign t[59] = ~(t[90] & t[91]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[92] | t[93]);
  assign t[61] = ~(t[211] | t[94]);
  assign t[62] = ~(t[95] ^ t[96]);
  assign t[63] = ~(t[97] | t[98]);
  assign t[64] = ~(t[212] | t[99]);
  assign t[65] = ~(t[100] ^ t[101]);
  assign t[66] = ~(t[213]);
  assign t[67] = ~(t[214]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[104] | t[105]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[215] | t[106]);
  assign t[71] = t[30] ? x[66] : x[65];
  assign t[72] = t[107] | t[52];
  assign t[73] = ~(t[108] | t[109]);
  assign t[74] = ~(t[216] | t[110]);
  assign t[75] = ~(t[111] | t[112]);
  assign t[76] = ~(t[113] ^ t[114]);
  assign t[77] = ~(t[115] | t[116]);
  assign t[78] = ~(t[217] | t[117]);
  assign t[79] = ~(t[118] | t[119]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[120] ^ t[121]);
  assign t[81] = ~(t[122]);
  assign t[82] = t[202] ? t[124] : t[123];
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = t[202] ? t[128] : t[127];
  assign t[85] = ~(t[218]);
  assign t[86] = ~(t[208] | t[209]);
  assign t[87] = ~(t[219]);
  assign t[88] = ~(t[220]);
  assign t[89] = ~(t[129] | t[130]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125] | t[131]);
  assign t[91] = ~(t[132]);
  assign t[92] = ~(t[221]);
  assign t[93] = ~(t[222]);
  assign t[94] = ~(t[133] | t[134]);
  assign t[95] = t[135] ? x[85] : x[84];
  assign t[96] = ~(t[136] & t[32]);
  assign t[97] = ~(t[223]);
  assign t[98] = ~(t[224]);
  assign t[99] = ~(t[137] | t[138]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [112:0] x;
 output y;

 wire [473:0] t;
  assign t[0] = t[1] ? t[2] : t[292];
  assign t[100] = ~(t[316]);
  assign t[101] = ~(t[317]);
  assign t[102] = ~(t[120] | t[121]);
  assign t[103] = ~(t[40]);
  assign t[104] = ~(t[122] | t[123]);
  assign t[105] = ~(t[124] & t[125]);
  assign t[106] = ~(t[318]);
  assign t[107] = ~(t[310] | t[311]);
  assign t[108] = ~(t[319]);
  assign t[109] = ~(t[320]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[126] | t[127]);
  assign t[111] = ~(t[114] | t[128]);
  assign t[112] = ~(t[321]);
  assign t[113] = ~(t[313] | t[314]);
  assign t[114] = ~(t[43] | t[129]);
  assign t[115] = ~(t[130]);
  assign t[116] = ~(t[131] & t[95]);
  assign t[117] = ~(t[132] & t[95]);
  assign t[118] = ~(t[97] & t[95]);
  assign t[119] = ~(t[294]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[322]);
  assign t[121] = ~(t[316] | t[317]);
  assign t[122] = ~(t[133] & t[42]);
  assign t[123] = t[29] | t[134];
  assign t[124] = t[296] & t[135];
  assign t[125] = t[131] | t[132];
  assign t[126] = ~(t[323]);
  assign t[127] = ~(t[319] | t[320]);
  assign t[128] = ~(t[136] & t[137]);
  assign t[129] = t[293] ? t[138] : t[116];
  assign t[12] = ~(t[18] ^ t[15]);
  assign t[130] = ~(t[139] | t[140]);
  assign t[131] = ~(x[7] | t[294]);
  assign t[132] = x[7] & t[294];
  assign t[133] = ~(t[135] & t[141]);
  assign t[134] = ~(t[43] | t[142]);
  assign t[135] = ~(t[67] | t[293]);
  assign t[136] = ~(t[143] | t[144]);
  assign t[137] = ~(t[67] & t[145]);
  assign t[138] = ~(t[132] & t[296]);
  assign t[139] = ~(t[43] | t[146]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = ~(t[43] | t[147]);
  assign t[141] = ~(t[69] & t[148]);
  assign t[142] = t[293] ? t[149] : t[117];
  assign t[143] = ~(t[67] | t[150]);
  assign t[144] = ~(t[43] | t[151]);
  assign t[145] = ~(t[68] & t[69]);
  assign t[146] = t[293] ? t[148] : t[118];
  assign t[147] = t[293] ? t[117] : t[149];
  assign t[148] = ~(x[7] & t[65]);
  assign t[149] = ~(t[131] & t[296]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[293] ? t[116] : t[117];
  assign t[151] = t[293] ? t[118] : t[148];
  assign t[152] = t[1] ? t[153] : t[298];
  assign t[153] = x[6] ? t[155] : t[154];
  assign t[154] = x[7] ? t[157] : t[156];
  assign t[155] = t[158] ^ x[86];
  assign t[156] = t[159] ^ t[160];
  assign t[157] = ~(t[161] ^ t[162]);
  assign t[158] = x[87] ^ x[88];
  assign t[159] = t[27] ? x[88] : x[87];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = ~(t[163] ^ t[162]);
  assign t[161] = x[7] ? t[165] : t[164];
  assign t[162] = ~(t[166] ^ t[167]);
  assign t[163] = x[7] ? t[169] : t[168];
  assign t[164] = ~(t[170] & t[171]);
  assign t[165] = t[159] ^ t[168];
  assign t[166] = x[7] ? t[173] : t[172];
  assign t[167] = x[7] ? t[175] : t[174];
  assign t[168] = ~(t[176] & t[177]);
  assign t[169] = t[178] ^ t[179];
  assign t[16] = ~(t[293] & t[294]);
  assign t[170] = ~(t[299] & t[46]);
  assign t[171] = ~(t[306] & t[180]);
  assign t[172] = ~(t[181] & t[182]);
  assign t[173] = t[183] ^ t[184];
  assign t[174] = ~(t[185] & t[186]);
  assign t[175] = t[187] ^ t[188];
  assign t[176] = ~(t[303] & t[57]);
  assign t[177] = ~(t[292] & t[189]);
  assign t[178] = t[27] ? x[90] : x[89];
  assign t[179] = ~(t[190] & t[191]);
  assign t[17] = ~(t[295] & t[296]);
  assign t[180] = ~(t[300] & t[45]);
  assign t[181] = ~(t[310] & t[80]);
  assign t[182] = ~(t[318] & t[192]);
  assign t[183] = t[103] ? x[92] : x[91];
  assign t[184] = ~(t[193] & t[194]);
  assign t[185] = ~(t[307] & t[73]);
  assign t[186] = ~(t[315] & t[195]);
  assign t[187] = t[103] ? x[94] : x[93];
  assign t[188] = ~(t[196] & t[197]);
  assign t[189] = ~(t[304] & t[56]);
  assign t[18] = x[7] ? t[26] : t[25];
  assign t[190] = ~(t[313] & t[89]);
  assign t[191] = ~(t[321] & t[198]);
  assign t[192] = ~(t[311] & t[79]);
  assign t[193] = ~(t[319] & t[109]);
  assign t[194] = ~(t[323] & t[199]);
  assign t[195] = ~(t[308] & t[72]);
  assign t[196] = ~(t[316] & t[101]);
  assign t[197] = ~(t[322] & t[200]);
  assign t[198] = ~(t[314] & t[88]);
  assign t[199] = ~(t[320] & t[108]);
  assign t[19] = t[27] ? x[10] : x[9];
  assign t[1] = ~(t[3]);
  assign t[200] = ~(t[317] & t[100]);
  assign t[201] = t[1] ? t[202] : t[303];
  assign t[202] = x[6] ? t[204] : t[203];
  assign t[203] = x[7] ? t[206] : t[205];
  assign t[204] = t[207] ^ x[95];
  assign t[205] = t[208] ^ t[209];
  assign t[206] = ~(t[210] ^ t[211]);
  assign t[207] = x[96] ^ x[97];
  assign t[208] = t[27] ? x[97] : x[96];
  assign t[209] = ~(t[212] ^ t[211]);
  assign t[20] = t[28] | t[29];
  assign t[210] = x[7] ? t[214] : t[213];
  assign t[211] = ~(t[215] ^ t[216]);
  assign t[212] = x[7] ? t[218] : t[217];
  assign t[213] = ~(t[219] & t[220]);
  assign t[214] = t[208] ^ t[217];
  assign t[215] = x[7] ? t[222] : t[221];
  assign t[216] = x[7] ? t[224] : t[223];
  assign t[217] = ~(t[225] & t[226]);
  assign t[218] = t[227] ^ t[228];
  assign t[219] = ~(t[46] & t[70]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[220] = ~(t[229] & t[297]);
  assign t[221] = ~(t[230] & t[231]);
  assign t[222] = t[232] ^ t[233];
  assign t[223] = ~(t[234] & t[235]);
  assign t[224] = t[236] ^ t[237];
  assign t[225] = ~(t[57] & t[86]);
  assign t[226] = ~(t[238] & t[298]);
  assign t[227] = t[27] ? x[99] : x[98];
  assign t[228] = ~(t[239] & t[240]);
  assign t[229] = ~(t[241] & t[45]);
  assign t[22] = ~(t[25] ^ t[13]);
  assign t[230] = ~(t[80] & t[106]);
  assign t[231] = ~(t[242] & t[302]);
  assign t[232] = t[103] ? x[101] : x[100];
  assign t[233] = ~(t[243] & t[244]);
  assign t[234] = ~(t[73] & t[98]);
  assign t[235] = ~(t[245] & t[301]);
  assign t[236] = t[103] ? x[103] : x[102];
  assign t[237] = ~(t[246] & t[247]);
  assign t[238] = ~(t[248] & t[56]);
  assign t[239] = ~(t[89] & t[112]);
  assign t[23] = x[7] ? t[33] : t[32];
  assign t[240] = ~(t[249] & t[305]);
  assign t[241] = ~(t[306] & t[300]);
  assign t[242] = ~(t[250] & t[79]);
  assign t[243] = ~(t[109] & t[126]);
  assign t[244] = ~(t[251] & t[312]);
  assign t[245] = ~(t[252] & t[72]);
  assign t[246] = ~(t[101] & t[120]);
  assign t[247] = ~(t[253] & t[309]);
  assign t[248] = ~(t[292] & t[304]);
  assign t[249] = ~(t[254] & t[88]);
  assign t[24] = x[7] ? t[35] : t[34];
  assign t[250] = ~(t[318] & t[311]);
  assign t[251] = ~(t[255] & t[108]);
  assign t[252] = ~(t[315] & t[308]);
  assign t[253] = ~(t[256] & t[100]);
  assign t[254] = ~(t[321] & t[314]);
  assign t[255] = ~(t[323] & t[320]);
  assign t[256] = ~(t[322] & t[317]);
  assign t[257] = t[1] ? t[258] : t[304];
  assign t[258] = x[6] ? t[260] : t[259];
  assign t[259] = x[7] ? t[262] : t[261];
  assign t[25] = ~(t[36] | t[37]);
  assign t[260] = t[263] ^ x[104];
  assign t[261] = t[264] ^ t[265];
  assign t[262] = ~(t[266] ^ t[267]);
  assign t[263] = x[105] ^ x[106];
  assign t[264] = t[27] ? x[106] : x[105];
  assign t[265] = ~(t[268] ^ t[267]);
  assign t[266] = x[7] ? t[270] : t[269];
  assign t[267] = ~(t[271] ^ t[272]);
  assign t[268] = x[7] ? t[274] : t[273];
  assign t[269] = ~(t[219] & t[275]);
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = t[264] ^ t[273];
  assign t[271] = x[7] ? t[277] : t[276];
  assign t[272] = x[7] ? t[279] : t[278];
  assign t[273] = ~(t[225] & t[280]);
  assign t[274] = t[281] ^ t[282];
  assign t[275] = t[30] | t[297];
  assign t[276] = ~(t[230] & t[283]);
  assign t[277] = t[284] ^ t[285];
  assign t[278] = ~(t[234] & t[286]);
  assign t[279] = t[287] ^ t[288];
  assign t[27] = ~(t[40]);
  assign t[280] = t[36] | t[298];
  assign t[281] = t[27] ? x[108] : x[107];
  assign t[282] = ~(t[239] & t[289]);
  assign t[283] = t[52] | t[302];
  assign t[284] = t[103] ? x[110] : x[109];
  assign t[285] = ~(t[243] & t[290]);
  assign t[286] = t[48] | t[301];
  assign t[287] = t[103] ? x[112] : x[111];
  assign t[288] = ~(t[246] & t[291]);
  assign t[289] = t[59] | t[305];
  assign t[28] = ~(t[41] & t[42]);
  assign t[290] = t[82] | t[312];
  assign t[291] = t[75] | t[309];
  assign t[292] = (t[324]);
  assign t[293] = (t[325]);
  assign t[294] = (t[326]);
  assign t[295] = (t[327]);
  assign t[296] = (t[328]);
  assign t[297] = (t[329]);
  assign t[298] = (t[330]);
  assign t[299] = (t[331]);
  assign t[29] = ~(t[43] | t[44]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (t[332]);
  assign t[301] = (t[333]);
  assign t[302] = (t[334]);
  assign t[303] = (t[335]);
  assign t[304] = (t[336]);
  assign t[305] = (t[337]);
  assign t[306] = (t[338]);
  assign t[307] = (t[339]);
  assign t[308] = (t[340]);
  assign t[309] = (t[341]);
  assign t[30] = ~(t[45] | t[46]);
  assign t[310] = (t[342]);
  assign t[311] = (t[343]);
  assign t[312] = (t[344]);
  assign t[313] = (t[345]);
  assign t[314] = (t[346]);
  assign t[315] = (t[347]);
  assign t[316] = (t[348]);
  assign t[317] = (t[349]);
  assign t[318] = (t[350]);
  assign t[319] = (t[351]);
  assign t[31] = ~(t[297] | t[47]);
  assign t[320] = (t[352]);
  assign t[321] = (t[353]);
  assign t[322] = (t[354]);
  assign t[323] = (t[355]);
  assign t[324] = t[356] ^ x[5];
  assign t[325] = t[357] ^ x[13];
  assign t[326] = t[358] ^ x[16];
  assign t[327] = t[359] ^ x[19];
  assign t[328] = t[360] ^ x[22];
  assign t[329] = t[361] ^ x[28];
  assign t[32] = ~(t[48] | t[49]);
  assign t[330] = t[362] ^ x[29];
  assign t[331] = t[363] ^ x[30];
  assign t[332] = t[364] ^ x[31];
  assign t[333] = t[365] ^ x[37];
  assign t[334] = t[366] ^ x[43];
  assign t[335] = t[367] ^ x[44];
  assign t[336] = t[368] ^ x[45];
  assign t[337] = t[369] ^ x[51];
  assign t[338] = t[370] ^ x[54];
  assign t[339] = t[371] ^ x[55];
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[340] = t[372] ^ x[56];
  assign t[341] = t[373] ^ x[62];
  assign t[342] = t[374] ^ x[65];
  assign t[343] = t[375] ^ x[66];
  assign t[344] = t[376] ^ x[72];
  assign t[345] = t[377] ^ x[75];
  assign t[346] = t[378] ^ x[76];
  assign t[347] = t[379] ^ x[77];
  assign t[348] = t[380] ^ x[78];
  assign t[349] = t[381] ^ x[79];
  assign t[34] = ~(t[52] | t[53]);
  assign t[350] = t[382] ^ x[80];
  assign t[351] = t[383] ^ x[81];
  assign t[352] = t[384] ^ x[82];
  assign t[353] = t[385] ^ x[83];
  assign t[354] = t[386] ^ x[84];
  assign t[355] = t[387] ^ x[85];
  assign t[356] = (~t[388] & t[389]);
  assign t[357] = (~t[390] & t[391]);
  assign t[358] = (~t[392] & t[393]);
  assign t[359] = (~t[394] & t[395]);
  assign t[35] = ~(t[54] ^ t[55]);
  assign t[360] = (~t[396] & t[397]);
  assign t[361] = (~t[398] & t[399]);
  assign t[362] = (~t[388] & t[400]);
  assign t[363] = (~t[398] & t[401]);
  assign t[364] = (~t[398] & t[402]);
  assign t[365] = (~t[403] & t[404]);
  assign t[366] = (~t[405] & t[406]);
  assign t[367] = (~t[388] & t[407]);
  assign t[368] = (~t[388] & t[408]);
  assign t[369] = (~t[409] & t[410]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[370] = (~t[398] & t[411]);
  assign t[371] = (~t[403] & t[412]);
  assign t[372] = (~t[403] & t[413]);
  assign t[373] = (~t[414] & t[415]);
  assign t[374] = (~t[405] & t[416]);
  assign t[375] = (~t[405] & t[417]);
  assign t[376] = (~t[418] & t[419]);
  assign t[377] = (~t[409] & t[420]);
  assign t[378] = (~t[409] & t[421]);
  assign t[379] = (~t[403] & t[422]);
  assign t[37] = ~(t[298] | t[58]);
  assign t[380] = (~t[414] & t[423]);
  assign t[381] = (~t[414] & t[424]);
  assign t[382] = (~t[405] & t[425]);
  assign t[383] = (~t[418] & t[426]);
  assign t[384] = (~t[418] & t[427]);
  assign t[385] = (~t[409] & t[428]);
  assign t[386] = (~t[414] & t[429]);
  assign t[387] = (~t[418] & t[430]);
  assign t[388] = t[431] ^ x[4];
  assign t[389] = t[432] ^ x[5];
  assign t[38] = ~(t[59] | t[60]);
  assign t[390] = t[433] ^ x[12];
  assign t[391] = t[434] ^ x[13];
  assign t[392] = t[435] ^ x[15];
  assign t[393] = t[436] ^ x[16];
  assign t[394] = t[437] ^ x[18];
  assign t[395] = t[438] ^ x[19];
  assign t[396] = t[439] ^ x[21];
  assign t[397] = t[440] ^ x[22];
  assign t[398] = t[441] ^ x[27];
  assign t[399] = t[442] ^ x[28];
  assign t[39] = ~(t[61] ^ t[62]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[443] ^ x[29];
  assign t[401] = t[444] ^ x[30];
  assign t[402] = t[445] ^ x[31];
  assign t[403] = t[446] ^ x[36];
  assign t[404] = t[447] ^ x[37];
  assign t[405] = t[448] ^ x[42];
  assign t[406] = t[449] ^ x[43];
  assign t[407] = t[450] ^ x[44];
  assign t[408] = t[451] ^ x[45];
  assign t[409] = t[452] ^ x[50];
  assign t[40] = ~(t[295]);
  assign t[410] = t[453] ^ x[51];
  assign t[411] = t[454] ^ x[54];
  assign t[412] = t[455] ^ x[55];
  assign t[413] = t[456] ^ x[56];
  assign t[414] = t[457] ^ x[61];
  assign t[415] = t[458] ^ x[62];
  assign t[416] = t[459] ^ x[65];
  assign t[417] = t[460] ^ x[66];
  assign t[418] = t[461] ^ x[71];
  assign t[419] = t[462] ^ x[72];
  assign t[41] = ~(t[63] | t[64]);
  assign t[420] = t[463] ^ x[75];
  assign t[421] = t[464] ^ x[76];
  assign t[422] = t[465] ^ x[77];
  assign t[423] = t[466] ^ x[78];
  assign t[424] = t[467] ^ x[79];
  assign t[425] = t[468] ^ x[80];
  assign t[426] = t[469] ^ x[81];
  assign t[427] = t[470] ^ x[82];
  assign t[428] = t[471] ^ x[83];
  assign t[429] = t[472] ^ x[84];
  assign t[42] = ~(t[65] & t[66]);
  assign t[430] = t[473] ^ x[85];
  assign t[431] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[432] = (x[0]);
  assign t[433] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[434] = (x[11]);
  assign t[435] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[436] = (x[14]);
  assign t[437] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[438] = (x[17]);
  assign t[439] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[43] = ~(t[67]);
  assign t[440] = (x[20]);
  assign t[441] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[442] = (x[24]);
  assign t[443] = (x[1]);
  assign t[444] = (x[25]);
  assign t[445] = (x[26]);
  assign t[446] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[447] = (x[33]);
  assign t[448] = (x[38] & ~x[39] & ~x[40] & ~x[41]) | (~x[38] & x[39] & ~x[40] & ~x[41]) | (~x[38] & ~x[39] & x[40] & ~x[41]) | (~x[38] & ~x[39] & ~x[40] & x[41]) | (x[38] & x[39] & x[40] & ~x[41]) | (x[38] & x[39] & ~x[40] & x[41]) | (x[38] & ~x[39] & x[40] & x[41]) | (~x[38] & x[39] & x[40] & x[41]);
  assign t[449] = (x[39]);
  assign t[44] = t[293] ? t[69] : t[68];
  assign t[450] = (x[2]);
  assign t[451] = (x[3]);
  assign t[452] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[453] = (x[47]);
  assign t[454] = (x[23]);
  assign t[455] = (x[34]);
  assign t[456] = (x[35]);
  assign t[457] = (x[57] & ~x[58] & ~x[59] & ~x[60]) | (~x[57] & x[58] & ~x[59] & ~x[60]) | (~x[57] & ~x[58] & x[59] & ~x[60]) | (~x[57] & ~x[58] & ~x[59] & x[60]) | (x[57] & x[58] & x[59] & ~x[60]) | (x[57] & x[58] & ~x[59] & x[60]) | (x[57] & ~x[58] & x[59] & x[60]) | (~x[57] & x[58] & x[59] & x[60]);
  assign t[458] = (x[58]);
  assign t[459] = (x[40]);
  assign t[45] = ~(t[299]);
  assign t[460] = (x[41]);
  assign t[461] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[462] = (x[68]);
  assign t[463] = (x[48]);
  assign t[464] = (x[49]);
  assign t[465] = (x[32]);
  assign t[466] = (x[59]);
  assign t[467] = (x[60]);
  assign t[468] = (x[38]);
  assign t[469] = (x[69]);
  assign t[46] = ~(t[300]);
  assign t[470] = (x[70]);
  assign t[471] = (x[46]);
  assign t[472] = (x[57]);
  assign t[473] = (x[67]);
  assign t[47] = ~(t[70] | t[71]);
  assign t[48] = ~(t[72] | t[73]);
  assign t[49] = ~(t[301] | t[74]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[75] | t[76]);
  assign t[51] = ~(t[77] ^ t[78]);
  assign t[52] = ~(t[79] | t[80]);
  assign t[53] = ~(t[302] | t[81]);
  assign t[54] = ~(t[82] | t[83]);
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = ~(t[303]);
  assign t[57] = ~(t[304]);
  assign t[58] = ~(t[86] | t[87]);
  assign t[59] = ~(t[88] | t[89]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[305] | t[90]);
  assign t[61] = t[27] ? x[53] : x[52];
  assign t[62] = ~(t[91] & t[92]);
  assign t[63] = ~(t[67] | t[93]);
  assign t[64] = ~(t[67] | t[94]);
  assign t[65] = ~(t[294] | t[95]);
  assign t[66] = t[43] & t[293];
  assign t[67] = ~(t[295]);
  assign t[68] = ~(x[7] & t[96]);
  assign t[69] = ~(t[296] & t[97]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[306]);
  assign t[71] = ~(t[299] | t[300]);
  assign t[72] = ~(t[307]);
  assign t[73] = ~(t[308]);
  assign t[74] = ~(t[98] | t[99]);
  assign t[75] = ~(t[100] | t[101]);
  assign t[76] = ~(t[309] | t[102]);
  assign t[77] = t[103] ? x[64] : x[63];
  assign t[78] = ~(t[104] & t[105]);
  assign t[79] = ~(t[310]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[311]);
  assign t[81] = ~(t[106] | t[107]);
  assign t[82] = ~(t[108] | t[109]);
  assign t[83] = ~(t[312] | t[110]);
  assign t[84] = t[103] ? x[74] : x[73];
  assign t[85] = ~(t[111] & t[42]);
  assign t[86] = ~(t[292]);
  assign t[87] = ~(t[303] | t[304]);
  assign t[88] = ~(t[313]);
  assign t[89] = ~(t[314]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[112] | t[113]);
  assign t[91] = ~(t[114]);
  assign t[92] = ~(t[115] | t[29]);
  assign t[93] = t[293] ? t[117] : t[116];
  assign t[94] = t[293] ? t[118] : t[68];
  assign t[95] = ~(t[296]);
  assign t[96] = ~(t[294] | t[296]);
  assign t[97] = ~(x[7] | t[119]);
  assign t[98] = ~(t[315]);
  assign t[99] = ~(t[307] | t[308]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[152] & ~t[201] & ~t[257]) | (~t[0] & t[152] & ~t[201] & ~t[257]) | (~t[0] & ~t[152] & t[201] & ~t[257]) | (~t[0] & ~t[152] & ~t[201] & t[257]) | (t[0] & t[152] & t[201] & ~t[257]) | (t[0] & t[152] & ~t[201] & t[257]) | (t[0] & ~t[152] & t[201] & t[257]) | (~t[0] & t[152] & t[201] & t[257]);
endmodule

module R2ind166(x, y);
 input [85:0] x;
 output y;

 wire [261:0] t;
  assign t[0] = t[1] ? t[2] : t[80];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = t[144] ^ x[5];
  assign t[113] = t[145] ^ x[13];
  assign t[114] = t[146] ^ x[16];
  assign t[115] = t[147] ^ x[19];
  assign t[116] = t[148] ^ x[22];
  assign t[117] = t[149] ^ x[28];
  assign t[118] = t[150] ^ x[29];
  assign t[119] = t[151] ^ x[32];
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[33];
  assign t[121] = t[153] ^ x[39];
  assign t[122] = t[154] ^ x[47];
  assign t[123] = t[155] ^ x[50];
  assign t[124] = t[156] ^ x[56];
  assign t[125] = t[157] ^ x[57];
  assign t[126] = t[158] ^ x[58];
  assign t[127] = t[159] ^ x[59];
  assign t[128] = t[160] ^ x[65];
  assign t[129] = t[161] ^ x[66];
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = t[162] ^ x[67];
  assign t[131] = t[163] ^ x[73];
  assign t[132] = t[164] ^ x[74];
  assign t[133] = t[165] ^ x[75];
  assign t[134] = t[166] ^ x[76];
  assign t[135] = t[167] ^ x[77];
  assign t[136] = t[168] ^ x[78];
  assign t[137] = t[169] ^ x[79];
  assign t[138] = t[170] ^ x[80];
  assign t[139] = t[171] ^ x[81];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[82];
  assign t[141] = t[173] ^ x[83];
  assign t[142] = t[174] ^ x[84];
  assign t[143] = t[175] ^ x[85];
  assign t[144] = (~t[176] & t[177]);
  assign t[145] = (~t[178] & t[179]);
  assign t[146] = (~t[180] & t[181]);
  assign t[147] = (~t[182] & t[183]);
  assign t[148] = (~t[184] & t[185]);
  assign t[149] = (~t[186] & t[187]);
  assign t[14] = x[7] ? t[21] : t[20];
  assign t[150] = (~t[176] & t[188]);
  assign t[151] = (~t[186] & t[189]);
  assign t[152] = (~t[186] & t[190]);
  assign t[153] = (~t[191] & t[192]);
  assign t[154] = (~t[193] & t[194]);
  assign t[155] = (~t[176] & t[195]);
  assign t[156] = (~t[196] & t[197]);
  assign t[157] = (~t[186] & t[198]);
  assign t[158] = (~t[191] & t[199]);
  assign t[159] = (~t[191] & t[200]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (~t[201] & t[202]);
  assign t[161] = (~t[193] & t[203]);
  assign t[162] = (~t[193] & t[204]);
  assign t[163] = (~t[205] & t[206]);
  assign t[164] = (~t[176] & t[207]);
  assign t[165] = (~t[196] & t[208]);
  assign t[166] = (~t[196] & t[209]);
  assign t[167] = (~t[191] & t[210]);
  assign t[168] = (~t[201] & t[211]);
  assign t[169] = (~t[201] & t[212]);
  assign t[16] = ~(t[81] & t[82]);
  assign t[170] = (~t[193] & t[213]);
  assign t[171] = (~t[205] & t[214]);
  assign t[172] = (~t[205] & t[215]);
  assign t[173] = (~t[196] & t[216]);
  assign t[174] = (~t[201] & t[217]);
  assign t[175] = (~t[205] & t[218]);
  assign t[176] = t[219] ^ x[4];
  assign t[177] = t[220] ^ x[5];
  assign t[178] = t[221] ^ x[12];
  assign t[179] = t[222] ^ x[13];
  assign t[17] = ~(t[83] & t[84]);
  assign t[180] = t[223] ^ x[15];
  assign t[181] = t[224] ^ x[16];
  assign t[182] = t[225] ^ x[18];
  assign t[183] = t[226] ^ x[19];
  assign t[184] = t[227] ^ x[21];
  assign t[185] = t[228] ^ x[22];
  assign t[186] = t[229] ^ x[27];
  assign t[187] = t[230] ^ x[28];
  assign t[188] = t[231] ^ x[29];
  assign t[189] = t[232] ^ x[32];
  assign t[18] = ~(t[24]);
  assign t[190] = t[233] ^ x[33];
  assign t[191] = t[234] ^ x[38];
  assign t[192] = t[235] ^ x[39];
  assign t[193] = t[236] ^ x[46];
  assign t[194] = t[237] ^ x[47];
  assign t[195] = t[238] ^ x[50];
  assign t[196] = t[239] ^ x[55];
  assign t[197] = t[240] ^ x[56];
  assign t[198] = t[241] ^ x[57];
  assign t[199] = t[242] ^ x[58];
  assign t[19] = x[7] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[59];
  assign t[201] = t[244] ^ x[64];
  assign t[202] = t[245] ^ x[65];
  assign t[203] = t[246] ^ x[66];
  assign t[204] = t[247] ^ x[67];
  assign t[205] = t[248] ^ x[72];
  assign t[206] = t[249] ^ x[73];
  assign t[207] = t[250] ^ x[74];
  assign t[208] = t[251] ^ x[75];
  assign t[209] = t[252] ^ x[76];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[253] ^ x[77];
  assign t[211] = t[254] ^ x[78];
  assign t[212] = t[255] ^ x[79];
  assign t[213] = t[256] ^ x[80];
  assign t[214] = t[257] ^ x[81];
  assign t[215] = t[258] ^ x[82];
  assign t[216] = t[259] ^ x[83];
  assign t[217] = t[260] ^ x[84];
  assign t[218] = t[261] ^ x[85];
  assign t[219] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[21] = t[12] ^ t[25];
  assign t[220] = (x[3]);
  assign t[221] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[222] = (x[11]);
  assign t[223] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[224] = (x[14]);
  assign t[225] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[226] = (x[17]);
  assign t[227] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[228] = (x[20]);
  assign t[229] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[22] = x[7] ? t[30] : t[29];
  assign t[230] = (x[24]);
  assign t[231] = (x[1]);
  assign t[232] = (x[26]);
  assign t[233] = (x[23]);
  assign t[234] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[235] = (x[35]);
  assign t[236] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[237] = (x[43]);
  assign t[238] = (x[0]);
  assign t[239] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[23] = x[7] ? t[32] : t[31];
  assign t[240] = (x[52]);
  assign t[241] = (x[25]);
  assign t[242] = (x[37]);
  assign t[243] = (x[34]);
  assign t[244] = (x[60] & ~x[61] & ~x[62] & ~x[63]) | (~x[60] & x[61] & ~x[62] & ~x[63]) | (~x[60] & ~x[61] & x[62] & ~x[63]) | (~x[60] & ~x[61] & ~x[62] & x[63]) | (x[60] & x[61] & x[62] & ~x[63]) | (x[60] & x[61] & ~x[62] & x[63]) | (x[60] & ~x[61] & x[62] & x[63]) | (~x[60] & x[61] & x[62] & x[63]);
  assign t[245] = (x[61]);
  assign t[246] = (x[45]);
  assign t[247] = (x[42]);
  assign t[248] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[249] = (x[69]);
  assign t[24] = ~(t[83]);
  assign t[250] = (x[2]);
  assign t[251] = (x[54]);
  assign t[252] = (x[51]);
  assign t[253] = (x[36]);
  assign t[254] = (x[63]);
  assign t[255] = (x[60]);
  assign t[256] = (x[44]);
  assign t[257] = (x[71]);
  assign t[258] = (x[68]);
  assign t[259] = (x[53]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[62]);
  assign t[261] = (x[70]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[37] & t[38]);
  assign t[28] = t[39] | t[85];
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] | t[86];
  assign t[35] = t[18] ? x[31] : x[30];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[87]);
  assign t[38] = ~(t[88]);
  assign t[39] = ~(t[53] | t[37]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[89];
  assign t[42] = t[57] ? x[41] : x[40];
  assign t[43] = ~(t[58] & t[59]);
  assign t[44] = ~(t[60] & t[61]);
  assign t[45] = t[62] | t[90];
  assign t[46] = t[57] ? x[49] : x[48];
  assign t[47] = ~(t[63] & t[64]);
  assign t[48] = ~(t[80]);
  assign t[49] = ~(t[91]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[65] | t[48]);
  assign t[51] = ~(t[66] & t[67]);
  assign t[52] = t[68] | t[92];
  assign t[53] = ~(t[93]);
  assign t[54] = ~(t[94]);
  assign t[55] = ~(t[95]);
  assign t[56] = ~(t[69] | t[54]);
  assign t[57] = ~(t[24]);
  assign t[58] = ~(t[70] & t[71]);
  assign t[59] = t[72] | t[96];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[97]);
  assign t[61] = ~(t[98]);
  assign t[62] = ~(t[73] | t[60]);
  assign t[63] = ~(t[74] & t[75]);
  assign t[64] = t[76] | t[99];
  assign t[65] = ~(t[100]);
  assign t[66] = ~(t[101]);
  assign t[67] = ~(t[102]);
  assign t[68] = ~(t[77] | t[66]);
  assign t[69] = ~(t[103]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104]);
  assign t[71] = ~(t[105]);
  assign t[72] = ~(t[78] | t[70]);
  assign t[73] = ~(t[106]);
  assign t[74] = ~(t[107]);
  assign t[75] = ~(t[108]);
  assign t[76] = ~(t[79] | t[74]);
  assign t[77] = ~(t[109]);
  assign t[78] = ~(t[110]);
  assign t[79] = ~(t[111]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[112]);
  assign t[81] = (t[113]);
  assign t[82] = (t[114]);
  assign t[83] = (t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [85:0] x;
 output y;

 wire [268:0] t;
  assign t[0] = t[1] ? t[2] : t[87];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = t[151] ^ x[5];
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[13];
  assign t[121] = t[153] ^ x[16];
  assign t[122] = t[154] ^ x[19];
  assign t[123] = t[155] ^ x[22];
  assign t[124] = t[156] ^ x[28];
  assign t[125] = t[157] ^ x[29];
  assign t[126] = t[158] ^ x[32];
  assign t[127] = t[159] ^ x[33];
  assign t[128] = t[160] ^ x[39];
  assign t[129] = t[161] ^ x[47];
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = t[162] ^ x[50];
  assign t[131] = t[163] ^ x[51];
  assign t[132] = t[164] ^ x[57];
  assign t[133] = t[165] ^ x[58];
  assign t[134] = t[166] ^ x[59];
  assign t[135] = t[167] ^ x[60];
  assign t[136] = t[168] ^ x[66];
  assign t[137] = t[169] ^ x[67];
  assign t[138] = t[170] ^ x[68];
  assign t[139] = t[171] ^ x[74];
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = t[172] ^ x[75];
  assign t[141] = t[173] ^ x[76];
  assign t[142] = t[174] ^ x[77];
  assign t[143] = t[175] ^ x[78];
  assign t[144] = t[176] ^ x[79];
  assign t[145] = t[177] ^ x[80];
  assign t[146] = t[178] ^ x[81];
  assign t[147] = t[179] ^ x[82];
  assign t[148] = t[180] ^ x[83];
  assign t[149] = t[181] ^ x[84];
  assign t[14] = x[7] ? t[21] : t[20];
  assign t[150] = t[182] ^ x[85];
  assign t[151] = (~t[183] & t[184]);
  assign t[152] = (~t[185] & t[186]);
  assign t[153] = (~t[187] & t[188]);
  assign t[154] = (~t[189] & t[190]);
  assign t[155] = (~t[191] & t[192]);
  assign t[156] = (~t[193] & t[194]);
  assign t[157] = (~t[183] & t[195]);
  assign t[158] = (~t[193] & t[196]);
  assign t[159] = (~t[193] & t[197]);
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = (~t[198] & t[199]);
  assign t[161] = (~t[200] & t[201]);
  assign t[162] = (~t[183] & t[202]);
  assign t[163] = (~t[183] & t[203]);
  assign t[164] = (~t[204] & t[205]);
  assign t[165] = (~t[193] & t[206]);
  assign t[166] = (~t[198] & t[207]);
  assign t[167] = (~t[198] & t[208]);
  assign t[168] = (~t[209] & t[210]);
  assign t[169] = (~t[200] & t[211]);
  assign t[16] = ~(t[88] & t[89]);
  assign t[170] = (~t[200] & t[212]);
  assign t[171] = (~t[213] & t[214]);
  assign t[172] = (~t[204] & t[215]);
  assign t[173] = (~t[204] & t[216]);
  assign t[174] = (~t[198] & t[217]);
  assign t[175] = (~t[209] & t[218]);
  assign t[176] = (~t[209] & t[219]);
  assign t[177] = (~t[200] & t[220]);
  assign t[178] = (~t[213] & t[221]);
  assign t[179] = (~t[213] & t[222]);
  assign t[17] = ~(t[90] & t[91]);
  assign t[180] = (~t[204] & t[223]);
  assign t[181] = (~t[209] & t[224]);
  assign t[182] = (~t[213] & t[225]);
  assign t[183] = t[226] ^ x[4];
  assign t[184] = t[227] ^ x[5];
  assign t[185] = t[228] ^ x[12];
  assign t[186] = t[229] ^ x[13];
  assign t[187] = t[230] ^ x[15];
  assign t[188] = t[231] ^ x[16];
  assign t[189] = t[232] ^ x[18];
  assign t[18] = ~(t[24]);
  assign t[190] = t[233] ^ x[19];
  assign t[191] = t[234] ^ x[21];
  assign t[192] = t[235] ^ x[22];
  assign t[193] = t[236] ^ x[27];
  assign t[194] = t[237] ^ x[28];
  assign t[195] = t[238] ^ x[29];
  assign t[196] = t[239] ^ x[32];
  assign t[197] = t[240] ^ x[33];
  assign t[198] = t[241] ^ x[38];
  assign t[199] = t[242] ^ x[39];
  assign t[19] = x[7] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[46];
  assign t[201] = t[244] ^ x[47];
  assign t[202] = t[245] ^ x[50];
  assign t[203] = t[246] ^ x[51];
  assign t[204] = t[247] ^ x[56];
  assign t[205] = t[248] ^ x[57];
  assign t[206] = t[249] ^ x[58];
  assign t[207] = t[250] ^ x[59];
  assign t[208] = t[251] ^ x[60];
  assign t[209] = t[252] ^ x[65];
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = t[253] ^ x[66];
  assign t[211] = t[254] ^ x[67];
  assign t[212] = t[255] ^ x[68];
  assign t[213] = t[256] ^ x[73];
  assign t[214] = t[257] ^ x[74];
  assign t[215] = t[258] ^ x[75];
  assign t[216] = t[259] ^ x[76];
  assign t[217] = t[260] ^ x[77];
  assign t[218] = t[261] ^ x[78];
  assign t[219] = t[262] ^ x[79];
  assign t[21] = t[12] ^ t[25];
  assign t[220] = t[263] ^ x[80];
  assign t[221] = t[264] ^ x[81];
  assign t[222] = t[265] ^ x[82];
  assign t[223] = t[266] ^ x[83];
  assign t[224] = t[267] ^ x[84];
  assign t[225] = t[268] ^ x[85];
  assign t[226] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[227] = (x[2]);
  assign t[228] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[229] = (x[11]);
  assign t[22] = x[7] ? t[30] : t[29];
  assign t[230] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[231] = (x[14]);
  assign t[232] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[233] = (x[17]);
  assign t[234] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[235] = (x[20]);
  assign t[236] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[237] = (x[24]);
  assign t[238] = (x[1]);
  assign t[239] = (x[26]);
  assign t[23] = x[7] ? t[32] : t[31];
  assign t[240] = (x[23]);
  assign t[241] = (x[34] & ~x[35] & ~x[36] & ~x[37]) | (~x[34] & x[35] & ~x[36] & ~x[37]) | (~x[34] & ~x[35] & x[36] & ~x[37]) | (~x[34] & ~x[35] & ~x[36] & x[37]) | (x[34] & x[35] & x[36] & ~x[37]) | (x[34] & x[35] & ~x[36] & x[37]) | (x[34] & ~x[35] & x[36] & x[37]) | (~x[34] & x[35] & x[36] & x[37]);
  assign t[242] = (x[35]);
  assign t[243] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[244] = (x[43]);
  assign t[245] = (x[3]);
  assign t[246] = (x[0]);
  assign t[247] = (x[52] & ~x[53] & ~x[54] & ~x[55]) | (~x[52] & x[53] & ~x[54] & ~x[55]) | (~x[52] & ~x[53] & x[54] & ~x[55]) | (~x[52] & ~x[53] & ~x[54] & x[55]) | (x[52] & x[53] & x[54] & ~x[55]) | (x[52] & x[53] & ~x[54] & x[55]) | (x[52] & ~x[53] & x[54] & x[55]) | (~x[52] & x[53] & x[54] & x[55]);
  assign t[248] = (x[53]);
  assign t[249] = (x[25]);
  assign t[24] = ~(t[90]);
  assign t[250] = (x[37]);
  assign t[251] = (x[34]);
  assign t[252] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[253] = (x[62]);
  assign t[254] = (x[45]);
  assign t[255] = (x[42]);
  assign t[256] = (x[69] & ~x[70] & ~x[71] & ~x[72]) | (~x[69] & x[70] & ~x[71] & ~x[72]) | (~x[69] & ~x[70] & x[71] & ~x[72]) | (~x[69] & ~x[70] & ~x[71] & x[72]) | (x[69] & x[70] & x[71] & ~x[72]) | (x[69] & x[70] & ~x[71] & x[72]) | (x[69] & ~x[70] & x[71] & x[72]) | (~x[69] & x[70] & x[71] & x[72]);
  assign t[257] = (x[70]);
  assign t[258] = (x[55]);
  assign t[259] = (x[52]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[260] = (x[36]);
  assign t[261] = (x[64]);
  assign t[262] = (x[61]);
  assign t[263] = (x[44]);
  assign t[264] = (x[72]);
  assign t[265] = (x[69]);
  assign t[266] = (x[54]);
  assign t[267] = (x[63]);
  assign t[268] = (x[71]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[37] & t[38]);
  assign t[28] = ~(t[39] & t[92]);
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = t[46] ^ t[47];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = ~(t[50] & t[93]);
  assign t[35] = t[18] ? x[31] : x[30];
  assign t[36] = ~(t[51] & t[52]);
  assign t[37] = ~(t[94]);
  assign t[38] = ~(t[95]);
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[55] & t[56]);
  assign t[41] = ~(t[57] & t[96]);
  assign t[42] = t[58] ? x[41] : x[40];
  assign t[43] = ~(t[59] & t[60]);
  assign t[44] = ~(t[61] & t[62]);
  assign t[45] = ~(t[63] & t[97]);
  assign t[46] = t[58] ? x[49] : x[48];
  assign t[47] = ~(t[64] & t[65]);
  assign t[48] = ~(t[98]);
  assign t[49] = ~(t[99]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[66] & t[67]);
  assign t[51] = ~(t[68] & t[69]);
  assign t[52] = ~(t[70] & t[100]);
  assign t[53] = ~(t[95] & t[94]);
  assign t[54] = ~(t[101]);
  assign t[55] = ~(t[102]);
  assign t[56] = ~(t[103]);
  assign t[57] = ~(t[71] & t[72]);
  assign t[58] = ~(t[24]);
  assign t[59] = ~(t[73] & t[74]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[75] & t[104]);
  assign t[61] = ~(t[105]);
  assign t[62] = ~(t[106]);
  assign t[63] = ~(t[76] & t[77]);
  assign t[64] = ~(t[78] & t[79]);
  assign t[65] = ~(t[80] & t[107]);
  assign t[66] = ~(t[99] & t[98]);
  assign t[67] = ~(t[87]);
  assign t[68] = ~(t[108]);
  assign t[69] = ~(t[109]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[81] & t[82]);
  assign t[71] = ~(t[103] & t[102]);
  assign t[72] = ~(t[110]);
  assign t[73] = ~(t[111]);
  assign t[74] = ~(t[112]);
  assign t[75] = ~(t[83] & t[84]);
  assign t[76] = ~(t[106] & t[105]);
  assign t[77] = ~(t[113]);
  assign t[78] = ~(t[114]);
  assign t[79] = ~(t[115]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[85] & t[86]);
  assign t[81] = ~(t[109] & t[108]);
  assign t[82] = ~(t[116]);
  assign t[83] = ~(t[112] & t[111]);
  assign t[84] = ~(t[117]);
  assign t[85] = ~(t[115] & t[114]);
  assign t[86] = ~(t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [79:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = t[1] ? t[2] : t[73];
  assign t[100] = t[126] ^ x[13];
  assign t[101] = t[127] ^ x[16];
  assign t[102] = t[128] ^ x[19];
  assign t[103] = t[129] ^ x[22];
  assign t[104] = t[130] ^ x[28];
  assign t[105] = t[131] ^ x[29];
  assign t[106] = t[132] ^ x[30];
  assign t[107] = t[133] ^ x[31];
  assign t[108] = t[134] ^ x[34];
  assign t[109] = t[135] ^ x[40];
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = t[136] ^ x[41];
  assign t[111] = t[137] ^ x[49];
  assign t[112] = t[138] ^ x[50];
  assign t[113] = t[139] ^ x[53];
  assign t[114] = t[140] ^ x[59];
  assign t[115] = t[141] ^ x[60];
  assign t[116] = t[142] ^ x[61];
  assign t[117] = t[143] ^ x[67];
  assign t[118] = t[144] ^ x[68];
  assign t[119] = t[145] ^ x[69];
  assign t[11] = ~(x[6]);
  assign t[120] = t[146] ^ x[75];
  assign t[121] = t[147] ^ x[76];
  assign t[122] = t[148] ^ x[77];
  assign t[123] = t[149] ^ x[78];
  assign t[124] = t[150] ^ x[79];
  assign t[125] = (~t[151] & t[152]);
  assign t[126] = (~t[153] & t[154]);
  assign t[127] = (~t[155] & t[156]);
  assign t[128] = (~t[157] & t[158]);
  assign t[129] = (~t[159] & t[160]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (~t[161] & t[162]);
  assign t[131] = (~t[161] & t[163]);
  assign t[132] = (~t[151] & t[164]);
  assign t[133] = (~t[151] & t[165]);
  assign t[134] = (~t[161] & t[166]);
  assign t[135] = (~t[167] & t[168]);
  assign t[136] = (~t[167] & t[169]);
  assign t[137] = (~t[170] & t[171]);
  assign t[138] = (~t[170] & t[172]);
  assign t[139] = (~t[151] & t[173]);
  assign t[13] = ~(t[19] ^ t[15]);
  assign t[140] = (~t[174] & t[175]);
  assign t[141] = (~t[174] & t[176]);
  assign t[142] = (~t[167] & t[177]);
  assign t[143] = (~t[178] & t[179]);
  assign t[144] = (~t[178] & t[180]);
  assign t[145] = (~t[170] & t[181]);
  assign t[146] = (~t[182] & t[183]);
  assign t[147] = (~t[182] & t[184]);
  assign t[148] = (~t[174] & t[185]);
  assign t[149] = (~t[178] & t[186]);
  assign t[14] = x[7] ? t[21] : t[20];
  assign t[150] = (~t[182] & t[187]);
  assign t[151] = t[188] ^ x[4];
  assign t[152] = t[189] ^ x[5];
  assign t[153] = t[190] ^ x[12];
  assign t[154] = t[191] ^ x[13];
  assign t[155] = t[192] ^ x[15];
  assign t[156] = t[193] ^ x[16];
  assign t[157] = t[194] ^ x[18];
  assign t[158] = t[195] ^ x[19];
  assign t[159] = t[196] ^ x[21];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[197] ^ x[22];
  assign t[161] = t[198] ^ x[27];
  assign t[162] = t[199] ^ x[28];
  assign t[163] = t[200] ^ x[29];
  assign t[164] = t[201] ^ x[30];
  assign t[165] = t[202] ^ x[31];
  assign t[166] = t[203] ^ x[34];
  assign t[167] = t[204] ^ x[39];
  assign t[168] = t[205] ^ x[40];
  assign t[169] = t[206] ^ x[41];
  assign t[16] = ~(t[74] & t[75]);
  assign t[170] = t[207] ^ x[48];
  assign t[171] = t[208] ^ x[49];
  assign t[172] = t[209] ^ x[50];
  assign t[173] = t[210] ^ x[53];
  assign t[174] = t[211] ^ x[58];
  assign t[175] = t[212] ^ x[59];
  assign t[176] = t[213] ^ x[60];
  assign t[177] = t[214] ^ x[61];
  assign t[178] = t[215] ^ x[66];
  assign t[179] = t[216] ^ x[67];
  assign t[17] = ~(t[76] & t[77]);
  assign t[180] = t[217] ^ x[68];
  assign t[181] = t[218] ^ x[69];
  assign t[182] = t[219] ^ x[74];
  assign t[183] = t[220] ^ x[75];
  assign t[184] = t[221] ^ x[76];
  assign t[185] = t[222] ^ x[77];
  assign t[186] = t[223] ^ x[78];
  assign t[187] = t[224] ^ x[79];
  assign t[188] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[189] = (x[1]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[191] = (x[11]);
  assign t[192] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[193] = (x[14]);
  assign t[194] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[195] = (x[17]);
  assign t[196] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[197] = (x[20]);
  assign t[198] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[199] = (x[25]);
  assign t[19] = x[7] ? t[26] : t[25];
  assign t[1] = ~(t[3]);
  assign t[200] = (x[23]);
  assign t[201] = (x[2]);
  assign t[202] = (x[0]);
  assign t[203] = (x[26]);
  assign t[204] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[205] = (x[37]);
  assign t[206] = (x[35]);
  assign t[207] = (x[44] & ~x[45] & ~x[46] & ~x[47]) | (~x[44] & x[45] & ~x[46] & ~x[47]) | (~x[44] & ~x[45] & x[46] & ~x[47]) | (~x[44] & ~x[45] & ~x[46] & x[47]) | (x[44] & x[45] & x[46] & ~x[47]) | (x[44] & x[45] & ~x[46] & x[47]) | (x[44] & ~x[45] & x[46] & x[47]) | (~x[44] & x[45] & x[46] & x[47]);
  assign t[208] = (x[46]);
  assign t[209] = (x[44]);
  assign t[20] = ~(t[27] & t[28]);
  assign t[210] = (x[3]);
  assign t[211] = (x[54] & ~x[55] & ~x[56] & ~x[57]) | (~x[54] & x[55] & ~x[56] & ~x[57]) | (~x[54] & ~x[55] & x[56] & ~x[57]) | (~x[54] & ~x[55] & ~x[56] & x[57]) | (x[54] & x[55] & x[56] & ~x[57]) | (x[54] & x[55] & ~x[56] & x[57]) | (x[54] & ~x[55] & x[56] & x[57]) | (~x[54] & x[55] & x[56] & x[57]);
  assign t[212] = (x[56]);
  assign t[213] = (x[54]);
  assign t[214] = (x[38]);
  assign t[215] = (x[62] & ~x[63] & ~x[64] & ~x[65]) | (~x[62] & x[63] & ~x[64] & ~x[65]) | (~x[62] & ~x[63] & x[64] & ~x[65]) | (~x[62] & ~x[63] & ~x[64] & x[65]) | (x[62] & x[63] & x[64] & ~x[65]) | (x[62] & x[63] & ~x[64] & x[65]) | (x[62] & ~x[63] & x[64] & x[65]) | (~x[62] & x[63] & x[64] & x[65]);
  assign t[216] = (x[64]);
  assign t[217] = (x[62]);
  assign t[218] = (x[47]);
  assign t[219] = (x[70] & ~x[71] & ~x[72] & ~x[73]) | (~x[70] & x[71] & ~x[72] & ~x[73]) | (~x[70] & ~x[71] & x[72] & ~x[73]) | (~x[70] & ~x[71] & ~x[72] & x[73]) | (x[70] & x[71] & x[72] & ~x[73]) | (x[70] & x[71] & ~x[72] & x[73]) | (x[70] & ~x[71] & x[72] & x[73]) | (~x[70] & x[71] & x[72] & x[73]);
  assign t[21] = t[12] ^ t[25];
  assign t[220] = (x[72]);
  assign t[221] = (x[70]);
  assign t[222] = (x[57]);
  assign t[223] = (x[65]);
  assign t[224] = (x[73]);
  assign t[22] = x[7] ? t[30] : t[29];
  assign t[23] = x[7] ? t[32] : t[31];
  assign t[24] = ~(t[76]);
  assign t[25] = ~(t[33] & t[34]);
  assign t[26] = t[35] ^ t[36];
  assign t[27] = ~(t[78] & t[37]);
  assign t[28] = ~(t[79] & t[38]);
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[43] & t[44]);
  assign t[32] = t[45] ^ t[46];
  assign t[33] = ~(t[80] & t[47]);
  assign t[34] = ~(t[81] & t[48]);
  assign t[35] = t[18] ? x[33] : x[32];
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = ~(t[82]);
  assign t[38] = ~(t[82] & t[51]);
  assign t[39] = ~(t[83] & t[52]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[84] & t[53]);
  assign t[41] = t[54] ? x[43] : x[42];
  assign t[42] = ~(t[55] & t[56]);
  assign t[43] = ~(t[85] & t[57]);
  assign t[44] = ~(t[86] & t[58]);
  assign t[45] = t[54] ? x[52] : x[51];
  assign t[46] = ~(t[59] & t[60]);
  assign t[47] = ~(t[87]);
  assign t[48] = ~(t[87] & t[61]);
  assign t[49] = ~(t[88] & t[62]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[89] & t[63]);
  assign t[51] = ~(t[78]);
  assign t[52] = ~(t[90]);
  assign t[53] = ~(t[90] & t[64]);
  assign t[54] = ~(t[24]);
  assign t[55] = ~(t[91] & t[65]);
  assign t[56] = ~(t[92] & t[66]);
  assign t[57] = ~(t[93]);
  assign t[58] = ~(t[93] & t[67]);
  assign t[59] = ~(t[94] & t[68]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[95] & t[69]);
  assign t[61] = ~(t[80]);
  assign t[62] = ~(t[96]);
  assign t[63] = ~(t[96] & t[70]);
  assign t[64] = ~(t[83]);
  assign t[65] = ~(t[97]);
  assign t[66] = ~(t[97] & t[71]);
  assign t[67] = ~(t[85]);
  assign t[68] = ~(t[98]);
  assign t[69] = ~(t[98] & t[72]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[88]);
  assign t[71] = ~(t[91]);
  assign t[72] = ~(t[94]);
  assign t[73] = (t[99]);
  assign t[74] = (t[100]);
  assign t[75] = (t[101]);
  assign t[76] = (t[102]);
  assign t[77] = (t[103]);
  assign t[78] = (t[104]);
  assign t[79] = (t[105]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[106]);
  assign t[81] = (t[107]);
  assign t[82] = (t[108]);
  assign t[83] = (t[109]);
  assign t[84] = (t[110]);
  assign t[85] = (t[111]);
  assign t[86] = (t[112]);
  assign t[87] = (t[113]);
  assign t[88] = (t[114]);
  assign t[89] = (t[115]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = (t[116]);
  assign t[91] = (t[117]);
  assign t[92] = (t[118]);
  assign t[93] = (t[119]);
  assign t[94] = (t[120]);
  assign t[95] = (t[121]);
  assign t[96] = (t[122]);
  assign t[97] = (t[123]);
  assign t[98] = (t[124]);
  assign t[99] = t[125] ^ x[5];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [85:0] x;
 output y;

 wire [333:0] t;
  assign t[0] = t[1] ? t[2] : t[152];
  assign t[100] = ~(t[176]);
  assign t[101] = ~(t[177]);
  assign t[102] = ~(t[120] | t[121]);
  assign t[103] = ~(t[40]);
  assign t[104] = ~(t[122] | t[123]);
  assign t[105] = ~(t[124] & t[125]);
  assign t[106] = ~(t[178]);
  assign t[107] = ~(t[170] | t[171]);
  assign t[108] = ~(t[179]);
  assign t[109] = ~(t[180]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[126] | t[127]);
  assign t[111] = ~(t[114] | t[128]);
  assign t[112] = ~(t[181]);
  assign t[113] = ~(t[173] | t[174]);
  assign t[114] = ~(t[43] | t[129]);
  assign t[115] = ~(t[130]);
  assign t[116] = ~(t[131] & t[95]);
  assign t[117] = ~(t[132] & t[95]);
  assign t[118] = ~(t[97] & t[95]);
  assign t[119] = ~(t[154]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[182]);
  assign t[121] = ~(t[176] | t[177]);
  assign t[122] = ~(t[133] & t[42]);
  assign t[123] = t[29] | t[134];
  assign t[124] = t[156] & t[135];
  assign t[125] = t[131] | t[132];
  assign t[126] = ~(t[183]);
  assign t[127] = ~(t[179] | t[180]);
  assign t[128] = ~(t[136] & t[137]);
  assign t[129] = t[153] ? t[138] : t[116];
  assign t[12] = ~(t[18] ^ t[15]);
  assign t[130] = ~(t[139] | t[140]);
  assign t[131] = ~(x[7] | t[154]);
  assign t[132] = x[7] & t[154];
  assign t[133] = ~(t[135] & t[141]);
  assign t[134] = ~(t[43] | t[142]);
  assign t[135] = ~(t[67] | t[153]);
  assign t[136] = ~(t[143] | t[144]);
  assign t[137] = ~(t[67] & t[145]);
  assign t[138] = ~(t[132] & t[156]);
  assign t[139] = ~(t[43] | t[146]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = ~(t[43] | t[147]);
  assign t[141] = ~(t[69] & t[148]);
  assign t[142] = t[153] ? t[149] : t[117];
  assign t[143] = ~(t[67] | t[150]);
  assign t[144] = ~(t[43] | t[151]);
  assign t[145] = ~(t[68] & t[69]);
  assign t[146] = t[153] ? t[148] : t[118];
  assign t[147] = t[153] ? t[117] : t[149];
  assign t[148] = ~(x[7] & t[65]);
  assign t[149] = ~(t[131] & t[156]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[153] ? t[116] : t[117];
  assign t[151] = t[153] ? t[118] : t[148];
  assign t[152] = (t[184]);
  assign t[153] = (t[185]);
  assign t[154] = (t[186]);
  assign t[155] = (t[187]);
  assign t[156] = (t[188]);
  assign t[157] = (t[189]);
  assign t[158] = (t[190]);
  assign t[159] = (t[191]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[192]);
  assign t[161] = (t[193]);
  assign t[162] = (t[194]);
  assign t[163] = (t[195]);
  assign t[164] = (t[196]);
  assign t[165] = (t[197]);
  assign t[166] = (t[198]);
  assign t[167] = (t[199]);
  assign t[168] = (t[200]);
  assign t[169] = (t[201]);
  assign t[16] = ~(t[153] & t[154]);
  assign t[170] = (t[202]);
  assign t[171] = (t[203]);
  assign t[172] = (t[204]);
  assign t[173] = (t[205]);
  assign t[174] = (t[206]);
  assign t[175] = (t[207]);
  assign t[176] = (t[208]);
  assign t[177] = (t[209]);
  assign t[178] = (t[210]);
  assign t[179] = (t[211]);
  assign t[17] = ~(t[155] & t[156]);
  assign t[180] = (t[212]);
  assign t[181] = (t[213]);
  assign t[182] = (t[214]);
  assign t[183] = (t[215]);
  assign t[184] = t[216] ^ x[5];
  assign t[185] = t[217] ^ x[13];
  assign t[186] = t[218] ^ x[16];
  assign t[187] = t[219] ^ x[19];
  assign t[188] = t[220] ^ x[22];
  assign t[189] = t[221] ^ x[28];
  assign t[18] = x[7] ? t[26] : t[25];
  assign t[190] = t[222] ^ x[29];
  assign t[191] = t[223] ^ x[30];
  assign t[192] = t[224] ^ x[31];
  assign t[193] = t[225] ^ x[37];
  assign t[194] = t[226] ^ x[43];
  assign t[195] = t[227] ^ x[44];
  assign t[196] = t[228] ^ x[45];
  assign t[197] = t[229] ^ x[51];
  assign t[198] = t[230] ^ x[54];
  assign t[199] = t[231] ^ x[55];
  assign t[19] = t[27] ? x[10] : x[9];
  assign t[1] = ~(t[3]);
  assign t[200] = t[232] ^ x[56];
  assign t[201] = t[233] ^ x[62];
  assign t[202] = t[234] ^ x[65];
  assign t[203] = t[235] ^ x[66];
  assign t[204] = t[236] ^ x[72];
  assign t[205] = t[237] ^ x[75];
  assign t[206] = t[238] ^ x[76];
  assign t[207] = t[239] ^ x[77];
  assign t[208] = t[240] ^ x[78];
  assign t[209] = t[241] ^ x[79];
  assign t[20] = t[28] | t[29];
  assign t[210] = t[242] ^ x[80];
  assign t[211] = t[243] ^ x[81];
  assign t[212] = t[244] ^ x[82];
  assign t[213] = t[245] ^ x[83];
  assign t[214] = t[246] ^ x[84];
  assign t[215] = t[247] ^ x[85];
  assign t[216] = (~t[248] & t[249]);
  assign t[217] = (~t[250] & t[251]);
  assign t[218] = (~t[252] & t[253]);
  assign t[219] = (~t[254] & t[255]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[220] = (~t[256] & t[257]);
  assign t[221] = (~t[258] & t[259]);
  assign t[222] = (~t[248] & t[260]);
  assign t[223] = (~t[258] & t[261]);
  assign t[224] = (~t[258] & t[262]);
  assign t[225] = (~t[263] & t[264]);
  assign t[226] = (~t[265] & t[266]);
  assign t[227] = (~t[248] & t[267]);
  assign t[228] = (~t[248] & t[268]);
  assign t[229] = (~t[269] & t[270]);
  assign t[22] = ~(t[25] ^ t[13]);
  assign t[230] = (~t[258] & t[271]);
  assign t[231] = (~t[263] & t[272]);
  assign t[232] = (~t[263] & t[273]);
  assign t[233] = (~t[274] & t[275]);
  assign t[234] = (~t[265] & t[276]);
  assign t[235] = (~t[265] & t[277]);
  assign t[236] = (~t[278] & t[279]);
  assign t[237] = (~t[269] & t[280]);
  assign t[238] = (~t[269] & t[281]);
  assign t[239] = (~t[263] & t[282]);
  assign t[23] = x[7] ? t[33] : t[32];
  assign t[240] = (~t[274] & t[283]);
  assign t[241] = (~t[274] & t[284]);
  assign t[242] = (~t[265] & t[285]);
  assign t[243] = (~t[278] & t[286]);
  assign t[244] = (~t[278] & t[287]);
  assign t[245] = (~t[269] & t[288]);
  assign t[246] = (~t[274] & t[289]);
  assign t[247] = (~t[278] & t[290]);
  assign t[248] = t[291] ^ x[4];
  assign t[249] = t[292] ^ x[5];
  assign t[24] = x[7] ? t[35] : t[34];
  assign t[250] = t[293] ^ x[12];
  assign t[251] = t[294] ^ x[13];
  assign t[252] = t[295] ^ x[15];
  assign t[253] = t[296] ^ x[16];
  assign t[254] = t[297] ^ x[18];
  assign t[255] = t[298] ^ x[19];
  assign t[256] = t[299] ^ x[21];
  assign t[257] = t[300] ^ x[22];
  assign t[258] = t[301] ^ x[27];
  assign t[259] = t[302] ^ x[28];
  assign t[25] = ~(t[36] | t[37]);
  assign t[260] = t[303] ^ x[29];
  assign t[261] = t[304] ^ x[30];
  assign t[262] = t[305] ^ x[31];
  assign t[263] = t[306] ^ x[36];
  assign t[264] = t[307] ^ x[37];
  assign t[265] = t[308] ^ x[42];
  assign t[266] = t[309] ^ x[43];
  assign t[267] = t[310] ^ x[44];
  assign t[268] = t[311] ^ x[45];
  assign t[269] = t[312] ^ x[50];
  assign t[26] = ~(t[38] ^ t[39]);
  assign t[270] = t[313] ^ x[51];
  assign t[271] = t[314] ^ x[54];
  assign t[272] = t[315] ^ x[55];
  assign t[273] = t[316] ^ x[56];
  assign t[274] = t[317] ^ x[61];
  assign t[275] = t[318] ^ x[62];
  assign t[276] = t[319] ^ x[65];
  assign t[277] = t[320] ^ x[66];
  assign t[278] = t[321] ^ x[71];
  assign t[279] = t[322] ^ x[72];
  assign t[27] = ~(t[40]);
  assign t[280] = t[323] ^ x[75];
  assign t[281] = t[324] ^ x[76];
  assign t[282] = t[325] ^ x[77];
  assign t[283] = t[326] ^ x[78];
  assign t[284] = t[327] ^ x[79];
  assign t[285] = t[328] ^ x[80];
  assign t[286] = t[329] ^ x[81];
  assign t[287] = t[330] ^ x[82];
  assign t[288] = t[331] ^ x[83];
  assign t[289] = t[332] ^ x[84];
  assign t[28] = ~(t[41] & t[42]);
  assign t[290] = t[333] ^ x[85];
  assign t[291] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[292] = (x[0]);
  assign t[293] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[294] = (x[11]);
  assign t[295] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[296] = (x[14]);
  assign t[297] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[298] = (x[17]);
  assign t[299] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[29] = ~(t[43] | t[44]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[20]);
  assign t[301] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[302] = (x[24]);
  assign t[303] = (x[1]);
  assign t[304] = (x[25]);
  assign t[305] = (x[26]);
  assign t[306] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[307] = (x[33]);
  assign t[308] = (x[38] & ~x[39] & ~x[40] & ~x[41]) | (~x[38] & x[39] & ~x[40] & ~x[41]) | (~x[38] & ~x[39] & x[40] & ~x[41]) | (~x[38] & ~x[39] & ~x[40] & x[41]) | (x[38] & x[39] & x[40] & ~x[41]) | (x[38] & x[39] & ~x[40] & x[41]) | (x[38] & ~x[39] & x[40] & x[41]) | (~x[38] & x[39] & x[40] & x[41]);
  assign t[309] = (x[39]);
  assign t[30] = ~(t[45] | t[46]);
  assign t[310] = (x[2]);
  assign t[311] = (x[3]);
  assign t[312] = (x[46] & ~x[47] & ~x[48] & ~x[49]) | (~x[46] & x[47] & ~x[48] & ~x[49]) | (~x[46] & ~x[47] & x[48] & ~x[49]) | (~x[46] & ~x[47] & ~x[48] & x[49]) | (x[46] & x[47] & x[48] & ~x[49]) | (x[46] & x[47] & ~x[48] & x[49]) | (x[46] & ~x[47] & x[48] & x[49]) | (~x[46] & x[47] & x[48] & x[49]);
  assign t[313] = (x[47]);
  assign t[314] = (x[23]);
  assign t[315] = (x[34]);
  assign t[316] = (x[35]);
  assign t[317] = (x[57] & ~x[58] & ~x[59] & ~x[60]) | (~x[57] & x[58] & ~x[59] & ~x[60]) | (~x[57] & ~x[58] & x[59] & ~x[60]) | (~x[57] & ~x[58] & ~x[59] & x[60]) | (x[57] & x[58] & x[59] & ~x[60]) | (x[57] & x[58] & ~x[59] & x[60]) | (x[57] & ~x[58] & x[59] & x[60]) | (~x[57] & x[58] & x[59] & x[60]);
  assign t[318] = (x[58]);
  assign t[319] = (x[40]);
  assign t[31] = ~(t[157] | t[47]);
  assign t[320] = (x[41]);
  assign t[321] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[322] = (x[68]);
  assign t[323] = (x[48]);
  assign t[324] = (x[49]);
  assign t[325] = (x[32]);
  assign t[326] = (x[59]);
  assign t[327] = (x[60]);
  assign t[328] = (x[38]);
  assign t[329] = (x[69]);
  assign t[32] = ~(t[48] | t[49]);
  assign t[330] = (x[70]);
  assign t[331] = (x[46]);
  assign t[332] = (x[57]);
  assign t[333] = (x[67]);
  assign t[33] = ~(t[50] ^ t[51]);
  assign t[34] = ~(t[52] | t[53]);
  assign t[35] = ~(t[54] ^ t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = ~(t[158] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = ~(t[61] ^ t[62]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[155]);
  assign t[41] = ~(t[63] | t[64]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = ~(t[67]);
  assign t[44] = t[153] ? t[69] : t[68];
  assign t[45] = ~(t[159]);
  assign t[46] = ~(t[160]);
  assign t[47] = ~(t[70] | t[71]);
  assign t[48] = ~(t[72] | t[73]);
  assign t[49] = ~(t[161] | t[74]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[75] | t[76]);
  assign t[51] = ~(t[77] ^ t[78]);
  assign t[52] = ~(t[79] | t[80]);
  assign t[53] = ~(t[162] | t[81]);
  assign t[54] = ~(t[82] | t[83]);
  assign t[55] = ~(t[84] ^ t[85]);
  assign t[56] = ~(t[163]);
  assign t[57] = ~(t[164]);
  assign t[58] = ~(t[86] | t[87]);
  assign t[59] = ~(t[88] | t[89]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[165] | t[90]);
  assign t[61] = t[27] ? x[53] : x[52];
  assign t[62] = ~(t[91] & t[92]);
  assign t[63] = ~(t[67] | t[93]);
  assign t[64] = ~(t[67] | t[94]);
  assign t[65] = ~(t[154] | t[95]);
  assign t[66] = t[43] & t[153];
  assign t[67] = ~(t[155]);
  assign t[68] = ~(x[7] & t[96]);
  assign t[69] = ~(t[156] & t[97]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[166]);
  assign t[71] = ~(t[159] | t[160]);
  assign t[72] = ~(t[167]);
  assign t[73] = ~(t[168]);
  assign t[74] = ~(t[98] | t[99]);
  assign t[75] = ~(t[100] | t[101]);
  assign t[76] = ~(t[169] | t[102]);
  assign t[77] = t[103] ? x[64] : x[63];
  assign t[78] = ~(t[104] & t[105]);
  assign t[79] = ~(t[170]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[171]);
  assign t[81] = ~(t[106] | t[107]);
  assign t[82] = ~(t[108] | t[109]);
  assign t[83] = ~(t[172] | t[110]);
  assign t[84] = t[103] ? x[74] : x[73];
  assign t[85] = ~(t[111] & t[42]);
  assign t[86] = ~(t[152]);
  assign t[87] = ~(t[163] | t[164]);
  assign t[88] = ~(t[173]);
  assign t[89] = ~(t[174]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[112] | t[113]);
  assign t[91] = ~(t[114]);
  assign t[92] = ~(t[115] | t[29]);
  assign t[93] = t[153] ? t[117] : t[116];
  assign t[94] = t[153] ? t[118] : t[68];
  assign t[95] = ~(t[156]);
  assign t[96] = ~(t[154] | t[156]);
  assign t[97] = ~(x[7] | t[119]);
  assign t[98] = ~(t[175]);
  assign t[99] = ~(t[167] | t[168]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [172:0] x;
 output y;

 wire [677:0] t;
  assign t[0] = t[1] ? t[2] : t[408];
  assign t[100] = ~(t[431]);
  assign t[101] = ~(t[144] | t[145]);
  assign t[102] = ~(t[146] | t[147]);
  assign t[103] = ~(t[432] | t[148]);
  assign t[104] = t[91] ? x[95] : x[94];
  assign t[105] = ~(t[149] & t[150]);
  assign t[106] = ~(t[433]);
  assign t[107] = ~(t[420] | t[421]);
  assign t[108] = ~(t[434]);
  assign t[109] = ~(t[435]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151] | t[152]);
  assign t[111] = ~(t[49]);
  assign t[112] = ~(t[137] | t[153]);
  assign t[113] = ~(t[154] | t[155]);
  assign t[114] = ~(t[436]);
  assign t[115] = ~(t[437]);
  assign t[116] = ~(t[156] | t[157]);
  assign t[117] = t[111] ? x[102] : x[101];
  assign t[118] = ~(t[158] & t[159]);
  assign t[119] = ~(t[438]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[439]);
  assign t[121] = ~(t[160] | t[161]);
  assign t[122] = ~(t[162] | t[163]);
  assign t[123] = ~(t[440] | t[164]);
  assign t[124] = t[111] ? x[112] : x[111];
  assign t[125] = ~(t[84] & t[149]);
  assign t[126] = ~(t[411]);
  assign t[127] = ~(t[165] & t[166]);
  assign t[128] = ~(x[7] & t[167]);
  assign t[129] = ~(t[81] | t[168]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[142] & t[169]);
  assign t[131] = ~(t[126] | t[170]);
  assign t[132] = ~(t[126] | t[171]);
  assign t[133] = ~(t[172] & t[412]);
  assign t[134] = ~(t[173] & t[166]);
  assign t[135] = ~(t[441]);
  assign t[136] = ~(t[426] | t[427]);
  assign t[137] = ~(t[81] | t[174]);
  assign t[138] = t[175] | t[176];
  assign t[139] = ~(t[177] & t[178]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[442]);
  assign t[141] = ~(t[428] | t[429]);
  assign t[142] = ~(t[179] | t[180]);
  assign t[143] = ~(t[181] | t[182]);
  assign t[144] = ~(t[443]);
  assign t[145] = ~(t[430] | t[431]);
  assign t[146] = ~(t[444]);
  assign t[147] = ~(t[445]);
  assign t[148] = ~(t[183] | t[184]);
  assign t[149] = ~(t[130] | t[185]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[129] | t[153]);
  assign t[151] = ~(t[446]);
  assign t[152] = ~(t[434] | t[435]);
  assign t[153] = ~(t[81] | t[186]);
  assign t[154] = t[412] & t[187];
  assign t[155] = ~(t[84]);
  assign t[156] = ~(t[447]);
  assign t[157] = ~(t[436] | t[437]);
  assign t[158] = ~(t[179] | t[132]);
  assign t[159] = ~(t[188] | t[176]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[448]);
  assign t[161] = ~(t[438] | t[439]);
  assign t[162] = ~(t[449]);
  assign t[163] = ~(t[450]);
  assign t[164] = ~(t[189] | t[190]);
  assign t[165] = ~(x[7] | t[191]);
  assign t[166] = ~(t[412]);
  assign t[167] = ~(t[410] | t[166]);
  assign t[168] = t[409] ? t[133] : t[134];
  assign t[169] = ~(t[126] & t[192]);
  assign t[16] = ~(t[409] & t[410]);
  assign t[170] = t[409] ? t[193] : t[134];
  assign t[171] = t[409] ? t[127] : t[194];
  assign t[172] = x[7] & t[410];
  assign t[173] = ~(x[7] | t[410]);
  assign t[174] = t[409] ? t[194] : t[195];
  assign t[175] = ~(t[84] & t[196]);
  assign t[176] = ~(t[81] | t[197]);
  assign t[177] = ~(t[198] | t[50]);
  assign t[178] = t[126] | t[199];
  assign t[179] = ~(t[126] | t[200]);
  assign t[17] = ~(t[411] & t[412]);
  assign t[180] = ~(t[81] | t[201]);
  assign t[181] = ~(t[81] | t[202]);
  assign t[182] = ~(t[150] & t[178]);
  assign t[183] = ~(t[451]);
  assign t[184] = ~(t[444] | t[445]);
  assign t[185] = ~(t[203] & t[178]);
  assign t[186] = t[409] ? t[193] : t[204];
  assign t[187] = ~(t[126] | t[409]);
  assign t[188] = ~(t[205]);
  assign t[189] = ~(t[452]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[449] | t[450]);
  assign t[191] = ~(t[410]);
  assign t[192] = ~(t[194] & t[195]);
  assign t[193] = ~(t[172] & t[166]);
  assign t[194] = ~(x[7] & t[206]);
  assign t[195] = ~(t[412] & t[165]);
  assign t[196] = ~(t[167] & t[207]);
  assign t[197] = t[409] ? t[195] : t[194];
  assign t[198] = ~(t[208]);
  assign t[199] = t[409] ? t[194] : t[127];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[409] ? t[134] : t[193];
  assign t[201] = t[409] ? t[127] : t[128];
  assign t[202] = t[409] ? t[204] : t[193];
  assign t[203] = ~(t[154] & t[209]);
  assign t[204] = ~(t[173] & t[412]);
  assign t[205] = ~(t[50] | t[153]);
  assign t[206] = ~(t[410] | t[412]);
  assign t[207] = t[81] & t[409];
  assign t[208] = ~(t[187] & t[210]);
  assign t[209] = t[173] | t[172];
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = ~(t[195] & t[128]);
  assign t[211] = t[1] ? t[212] : t[453];
  assign t[212] = x[6] ? t[214] : t[213];
  assign t[213] = x[7] ? t[216] : t[215];
  assign t[214] = t[217] ^ x[126];
  assign t[215] = t[218] ^ t[219];
  assign t[216] = ~(t[220] ^ t[221]);
  assign t[217] = x[127] ^ x[128];
  assign t[218] = t[30] ? x[128] : x[127];
  assign t[219] = ~(t[222] ^ t[223]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = x[7] ? t[225] : t[224];
  assign t[221] = ~(t[226] ^ t[227]);
  assign t[222] = x[7] ? t[229] : t[228];
  assign t[223] = ~(t[230] ^ t[231]);
  assign t[224] = ~(t[232] & t[233]);
  assign t[225] = t[234] ^ t[235];
  assign t[226] = x[7] ? t[237] : t[236];
  assign t[227] = x[7] ? t[239] : t[238];
  assign t[228] = ~(t[240] & t[241]);
  assign t[229] = t[242] ^ t[243];
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = x[7] ? t[245] : t[244];
  assign t[231] = x[7] ? t[247] : t[246];
  assign t[232] = ~(t[415] & t[54]);
  assign t[233] = ~(t[425] & t[248]);
  assign t[234] = t[91] ? x[130] : x[129];
  assign t[235] = ~(t[249] & t[250]);
  assign t[236] = ~(t[251] & t[252]);
  assign t[237] = t[253] ^ t[254];
  assign t[238] = ~(t[255] & t[256]);
  assign t[239] = t[257] ^ t[244];
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = ~(t[420] & t[68]);
  assign t[241] = ~(t[433] & t[258]);
  assign t[242] = t[111] ? x[132] : x[131];
  assign t[243] = ~(t[259] & t[260]);
  assign t[244] = ~(t[261] & t[262]);
  assign t[245] = t[263] ^ t[264];
  assign t[246] = ~(t[265] & t[266]);
  assign t[247] = t[267] ^ t[246];
  assign t[248] = ~(t[416] & t[53]);
  assign t[249] = ~(t[426] & t[89]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = ~(t[441] & t[268]);
  assign t[251] = ~(t[430] & t[100]);
  assign t[252] = ~(t[443] & t[269]);
  assign t[253] = t[111] ? x[134] : x[133];
  assign t[254] = ~(t[270] & t[271]);
  assign t[255] = ~(t[428] & t[95]);
  assign t[256] = ~(t[442] & t[272]);
  assign t[257] = t[91] ? x[136] : x[135];
  assign t[258] = ~(t[421] & t[67]);
  assign t[259] = ~(t[434] & t[109]);
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = ~(t[446] & t[273]);
  assign t[261] = ~(t[438] & t[120]);
  assign t[262] = ~(t[448] & t[274]);
  assign t[263] = t[111] ? x[138] : x[137];
  assign t[264] = ~(t[275] & t[276]);
  assign t[265] = ~(t[436] & t[115]);
  assign t[266] = ~(t[447] & t[277]);
  assign t[267] = t[111] ? x[140] : x[139];
  assign t[268] = ~(t[427] & t[88]);
  assign t[269] = ~(t[431] & t[99]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = ~(t[444] & t[147]);
  assign t[271] = ~(t[451] & t[278]);
  assign t[272] = ~(t[429] & t[94]);
  assign t[273] = ~(t[435] & t[108]);
  assign t[274] = ~(t[439] & t[119]);
  assign t[275] = ~(t[449] & t[163]);
  assign t[276] = ~(t[452] & t[279]);
  assign t[277] = ~(t[437] & t[114]);
  assign t[278] = ~(t[445] & t[146]);
  assign t[279] = ~(t[450] & t[162]);
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[1] ? t[281] : t[454];
  assign t[281] = x[6] ? t[283] : t[282];
  assign t[282] = x[7] ? t[285] : t[284];
  assign t[283] = t[286] ^ x[142];
  assign t[284] = t[287] ^ t[288];
  assign t[285] = ~(t[289] ^ t[290]);
  assign t[286] = x[143] ^ x[144];
  assign t[287] = t[30] ? x[144] : x[143];
  assign t[288] = ~(t[291] ^ t[292]);
  assign t[289] = x[7] ? t[294] : t[293];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = ~(t[295] ^ t[296]);
  assign t[291] = x[7] ? t[298] : t[297];
  assign t[292] = ~(t[299] ^ t[300]);
  assign t[293] = ~(t[301] & t[302]);
  assign t[294] = t[303] ^ t[304];
  assign t[295] = x[7] ? t[306] : t[305];
  assign t[296] = x[7] ? t[308] : t[307];
  assign t[297] = ~(t[309] & t[310]);
  assign t[298] = t[311] ^ t[312];
  assign t[299] = x[7] ? t[314] : t[313];
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = x[7] ? t[316] : t[315];
  assign t[301] = ~(t[54] & t[86]);
  assign t[302] = ~(t[317] & t[413]);
  assign t[303] = t[91] ? x[146] : x[145];
  assign t[304] = ~(t[318] & t[319]);
  assign t[305] = ~(t[320] & t[321]);
  assign t[306] = t[322] ^ t[323];
  assign t[307] = ~(t[324] & t[325]);
  assign t[308] = t[326] ^ t[315];
  assign t[309] = ~(t[68] & t[106]);
  assign t[30] = ~(t[49]);
  assign t[310] = ~(t[327] & t[414]);
  assign t[311] = t[111] ? x[148] : x[147];
  assign t[312] = ~(t[328] & t[329]);
  assign t[313] = ~(t[330] & t[331]);
  assign t[314] = t[332] ^ t[313];
  assign t[315] = ~(t[333] & t[334]);
  assign t[316] = t[335] ^ t[336];
  assign t[317] = ~(t[337] & t[53]);
  assign t[318] = ~(t[89] & t[135]);
  assign t[319] = ~(t[338] & t[417]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = ~(t[100] & t[144]);
  assign t[321] = ~(t[339] & t[419]);
  assign t[322] = t[91] ? x[150] : x[149];
  assign t[323] = ~(t[340] & t[341]);
  assign t[324] = ~(t[95] & t[140]);
  assign t[325] = ~(t[342] & t[418]);
  assign t[326] = t[30] ? x[152] : x[151];
  assign t[327] = ~(t[343] & t[67]);
  assign t[328] = ~(t[109] & t[151]);
  assign t[329] = ~(t[344] & t[422]);
  assign t[32] = ~(t[52]);
  assign t[330] = ~(t[115] & t[156]);
  assign t[331] = ~(t[345] & t[423]);
  assign t[332] = t[111] ? x[154] : x[153];
  assign t[333] = ~(t[120] & t[160]);
  assign t[334] = ~(t[346] & t[424]);
  assign t[335] = t[111] ? x[156] : x[155];
  assign t[336] = ~(t[347] & t[348]);
  assign t[337] = ~(t[425] & t[416]);
  assign t[338] = ~(t[349] & t[88]);
  assign t[339] = ~(t[350] & t[99]);
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = ~(t[147] & t[183]);
  assign t[341] = ~(t[351] & t[432]);
  assign t[342] = ~(t[352] & t[94]);
  assign t[343] = ~(t[433] & t[421]);
  assign t[344] = ~(t[353] & t[108]);
  assign t[345] = ~(t[354] & t[114]);
  assign t[346] = ~(t[355] & t[119]);
  assign t[347] = ~(t[163] & t[189]);
  assign t[348] = ~(t[356] & t[440]);
  assign t[349] = ~(t[441] & t[427]);
  assign t[34] = ~(t[413] | t[55]);
  assign t[350] = ~(t[443] & t[431]);
  assign t[351] = ~(t[357] & t[146]);
  assign t[352] = ~(t[442] & t[429]);
  assign t[353] = ~(t[446] & t[435]);
  assign t[354] = ~(t[447] & t[437]);
  assign t[355] = ~(t[448] & t[439]);
  assign t[356] = ~(t[358] & t[162]);
  assign t[357] = ~(t[451] & t[445]);
  assign t[358] = ~(t[452] & t[450]);
  assign t[359] = t[1] ? t[360] : t[455];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = x[6] ? t[362] : t[361];
  assign t[361] = x[7] ? t[364] : t[363];
  assign t[362] = t[365] ^ x[158];
  assign t[363] = t[366] ^ t[367];
  assign t[364] = ~(t[368] ^ t[369]);
  assign t[365] = x[159] ^ x[160];
  assign t[366] = t[30] ? x[160] : x[159];
  assign t[367] = ~(t[370] ^ t[371]);
  assign t[368] = x[7] ? t[373] : t[372];
  assign t[369] = ~(t[374] ^ t[375]);
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = x[7] ? t[377] : t[376];
  assign t[371] = ~(t[378] ^ t[379]);
  assign t[372] = ~(t[301] & t[380]);
  assign t[373] = t[381] ^ t[382];
  assign t[374] = x[7] ? t[384] : t[383];
  assign t[375] = x[7] ? t[386] : t[385];
  assign t[376] = ~(t[309] & t[387]);
  assign t[377] = t[388] ^ t[389];
  assign t[378] = x[7] ? t[391] : t[390];
  assign t[379] = x[7] ? t[393] : t[392];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[33] | t[413];
  assign t[381] = t[91] ? x[162] : x[161];
  assign t[382] = ~(t[318] & t[394]);
  assign t[383] = ~(t[320] & t[395]);
  assign t[384] = t[396] ^ t[397];
  assign t[385] = ~(t[324] & t[398]);
  assign t[386] = t[399] ^ t[392];
  assign t[387] = t[41] | t[414];
  assign t[388] = t[111] ? x[164] : x[163];
  assign t[389] = ~(t[328] & t[400]);
  assign t[38] = ~(t[47] ^ t[62]);
  assign t[390] = ~(t[330] & t[401]);
  assign t[391] = t[402] ^ t[390];
  assign t[392] = ~(t[333] & t[403]);
  assign t[393] = t[404] ^ t[405];
  assign t[394] = t[56] | t[417];
  assign t[395] = t[63] | t[419];
  assign t[396] = t[91] ? x[166] : x[165];
  assign t[397] = ~(t[340] & t[406]);
  assign t[398] = t[60] | t[418];
  assign t[399] = t[111] ? x[168] : x[167];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[70] | t[422];
  assign t[401] = t[74] | t[423];
  assign t[402] = t[111] ? x[170] : x[169];
  assign t[403] = t[77] | t[424];
  assign t[404] = t[111] ? x[172] : x[171];
  assign t[405] = ~(t[347] & t[407]);
  assign t[406] = t[102] | t[432];
  assign t[407] = t[122] | t[440];
  assign t[408] = (t[456]);
  assign t[409] = (t[457]);
  assign t[40] = ~(t[65] ^ t[66]);
  assign t[410] = (t[458]);
  assign t[411] = (t[459]);
  assign t[412] = (t[460]);
  assign t[413] = (t[461]);
  assign t[414] = (t[462]);
  assign t[415] = (t[463]);
  assign t[416] = (t[464]);
  assign t[417] = (t[465]);
  assign t[418] = (t[466]);
  assign t[419] = (t[467]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[420] = (t[468]);
  assign t[421] = (t[469]);
  assign t[422] = (t[470]);
  assign t[423] = (t[471]);
  assign t[424] = (t[472]);
  assign t[425] = (t[473]);
  assign t[426] = (t[474]);
  assign t[427] = (t[475]);
  assign t[428] = (t[476]);
  assign t[429] = (t[477]);
  assign t[42] = ~(t[414] | t[69]);
  assign t[430] = (t[478]);
  assign t[431] = (t[479]);
  assign t[432] = (t[480]);
  assign t[433] = (t[481]);
  assign t[434] = (t[482]);
  assign t[435] = (t[483]);
  assign t[436] = (t[484]);
  assign t[437] = (t[485]);
  assign t[438] = (t[486]);
  assign t[439] = (t[487]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (t[488]);
  assign t[441] = (t[489]);
  assign t[442] = (t[490]);
  assign t[443] = (t[491]);
  assign t[444] = (t[492]);
  assign t[445] = (t[493]);
  assign t[446] = (t[494]);
  assign t[447] = (t[495]);
  assign t[448] = (t[496]);
  assign t[449] = (t[497]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (t[498]);
  assign t[451] = (t[499]);
  assign t[452] = (t[500]);
  assign t[453] = (t[501]);
  assign t[454] = (t[502]);
  assign t[455] = (t[503]);
  assign t[456] = t[504] ^ x[5];
  assign t[457] = t[505] ^ x[13];
  assign t[458] = t[506] ^ x[16];
  assign t[459] = t[507] ^ x[19];
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = t[508] ^ x[22];
  assign t[461] = t[509] ^ x[28];
  assign t[462] = t[510] ^ x[34];
  assign t[463] = t[511] ^ x[35];
  assign t[464] = t[512] ^ x[36];
  assign t[465] = t[513] ^ x[42];
  assign t[466] = t[514] ^ x[50];
  assign t[467] = t[515] ^ x[56];
  assign t[468] = t[516] ^ x[57];
  assign t[469] = t[517] ^ x[58];
  assign t[46] = ~(t[45] ^ t[76]);
  assign t[470] = t[518] ^ x[64];
  assign t[471] = t[519] ^ x[72];
  assign t[472] = t[520] ^ x[78];
  assign t[473] = t[521] ^ x[79];
  assign t[474] = t[522] ^ x[80];
  assign t[475] = t[523] ^ x[81];
  assign t[476] = t[524] ^ x[82];
  assign t[477] = t[525] ^ x[83];
  assign t[478] = t[526] ^ x[86];
  assign t[479] = t[527] ^ x[87];
  assign t[47] = ~(t[77] | t[78]);
  assign t[480] = t[528] ^ x[93];
  assign t[481] = t[529] ^ x[96];
  assign t[482] = t[530] ^ x[97];
  assign t[483] = t[531] ^ x[98];
  assign t[484] = t[532] ^ x[99];
  assign t[485] = t[533] ^ x[100];
  assign t[486] = t[534] ^ x[103];
  assign t[487] = t[535] ^ x[104];
  assign t[488] = t[536] ^ x[110];
  assign t[489] = t[537] ^ x[113];
  assign t[48] = ~(t[79] ^ t[80]);
  assign t[490] = t[538] ^ x[114];
  assign t[491] = t[539] ^ x[115];
  assign t[492] = t[540] ^ x[116];
  assign t[493] = t[541] ^ x[117];
  assign t[494] = t[542] ^ x[118];
  assign t[495] = t[543] ^ x[119];
  assign t[496] = t[544] ^ x[120];
  assign t[497] = t[545] ^ x[121];
  assign t[498] = t[546] ^ x[122];
  assign t[499] = t[547] ^ x[123];
  assign t[49] = ~(t[411]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = t[548] ^ x[124];
  assign t[501] = t[549] ^ x[125];
  assign t[502] = t[550] ^ x[141];
  assign t[503] = t[551] ^ x[157];
  assign t[504] = (~t[552] & t[553]);
  assign t[505] = (~t[554] & t[555]);
  assign t[506] = (~t[556] & t[557]);
  assign t[507] = (~t[558] & t[559]);
  assign t[508] = (~t[560] & t[561]);
  assign t[509] = (~t[562] & t[563]);
  assign t[50] = ~(t[81] | t[82]);
  assign t[510] = (~t[564] & t[565]);
  assign t[511] = (~t[562] & t[566]);
  assign t[512] = (~t[562] & t[567]);
  assign t[513] = (~t[568] & t[569]);
  assign t[514] = (~t[570] & t[571]);
  assign t[515] = (~t[572] & t[573]);
  assign t[516] = (~t[564] & t[574]);
  assign t[517] = (~t[564] & t[575]);
  assign t[518] = (~t[576] & t[577]);
  assign t[519] = (~t[578] & t[579]);
  assign t[51] = ~(t[83] & t[84]);
  assign t[520] = (~t[580] & t[581]);
  assign t[521] = (~t[562] & t[582]);
  assign t[522] = (~t[568] & t[583]);
  assign t[523] = (~t[568] & t[584]);
  assign t[524] = (~t[570] & t[585]);
  assign t[525] = (~t[570] & t[586]);
  assign t[526] = (~t[572] & t[587]);
  assign t[527] = (~t[572] & t[588]);
  assign t[528] = (~t[589] & t[590]);
  assign t[529] = (~t[564] & t[591]);
  assign t[52] = ~(t[81] | t[85]);
  assign t[530] = (~t[576] & t[592]);
  assign t[531] = (~t[576] & t[593]);
  assign t[532] = (~t[578] & t[594]);
  assign t[533] = (~t[578] & t[595]);
  assign t[534] = (~t[580] & t[596]);
  assign t[535] = (~t[580] & t[597]);
  assign t[536] = (~t[598] & t[599]);
  assign t[537] = (~t[568] & t[600]);
  assign t[538] = (~t[570] & t[601]);
  assign t[539] = (~t[572] & t[602]);
  assign t[53] = ~(t[415]);
  assign t[540] = (~t[589] & t[603]);
  assign t[541] = (~t[589] & t[604]);
  assign t[542] = (~t[576] & t[605]);
  assign t[543] = (~t[578] & t[606]);
  assign t[544] = (~t[580] & t[607]);
  assign t[545] = (~t[598] & t[608]);
  assign t[546] = (~t[598] & t[609]);
  assign t[547] = (~t[589] & t[610]);
  assign t[548] = (~t[598] & t[611]);
  assign t[549] = (~t[552] & t[612]);
  assign t[54] = ~(t[416]);
  assign t[550] = (~t[552] & t[613]);
  assign t[551] = (~t[552] & t[614]);
  assign t[552] = t[615] ^ x[4];
  assign t[553] = t[616] ^ x[5];
  assign t[554] = t[617] ^ x[12];
  assign t[555] = t[618] ^ x[13];
  assign t[556] = t[619] ^ x[15];
  assign t[557] = t[620] ^ x[16];
  assign t[558] = t[621] ^ x[18];
  assign t[559] = t[622] ^ x[19];
  assign t[55] = ~(t[86] | t[87]);
  assign t[560] = t[623] ^ x[21];
  assign t[561] = t[624] ^ x[22];
  assign t[562] = t[625] ^ x[27];
  assign t[563] = t[626] ^ x[28];
  assign t[564] = t[627] ^ x[33];
  assign t[565] = t[628] ^ x[34];
  assign t[566] = t[629] ^ x[35];
  assign t[567] = t[630] ^ x[36];
  assign t[568] = t[631] ^ x[41];
  assign t[569] = t[632] ^ x[42];
  assign t[56] = ~(t[88] | t[89]);
  assign t[570] = t[633] ^ x[49];
  assign t[571] = t[634] ^ x[50];
  assign t[572] = t[635] ^ x[55];
  assign t[573] = t[636] ^ x[56];
  assign t[574] = t[637] ^ x[57];
  assign t[575] = t[638] ^ x[58];
  assign t[576] = t[639] ^ x[63];
  assign t[577] = t[640] ^ x[64];
  assign t[578] = t[641] ^ x[71];
  assign t[579] = t[642] ^ x[72];
  assign t[57] = ~(t[417] | t[90]);
  assign t[580] = t[643] ^ x[77];
  assign t[581] = t[644] ^ x[78];
  assign t[582] = t[645] ^ x[79];
  assign t[583] = t[646] ^ x[80];
  assign t[584] = t[647] ^ x[81];
  assign t[585] = t[648] ^ x[82];
  assign t[586] = t[649] ^ x[83];
  assign t[587] = t[650] ^ x[86];
  assign t[588] = t[651] ^ x[87];
  assign t[589] = t[652] ^ x[92];
  assign t[58] = t[91] ? x[44] : x[43];
  assign t[590] = t[653] ^ x[93];
  assign t[591] = t[654] ^ x[96];
  assign t[592] = t[655] ^ x[97];
  assign t[593] = t[656] ^ x[98];
  assign t[594] = t[657] ^ x[99];
  assign t[595] = t[658] ^ x[100];
  assign t[596] = t[659] ^ x[103];
  assign t[597] = t[660] ^ x[104];
  assign t[598] = t[661] ^ x[109];
  assign t[599] = t[662] ^ x[110];
  assign t[59] = ~(t[92] & t[93]);
  assign t[5] = t[9] ^ x[8];
  assign t[600] = t[663] ^ x[113];
  assign t[601] = t[664] ^ x[114];
  assign t[602] = t[665] ^ x[115];
  assign t[603] = t[666] ^ x[116];
  assign t[604] = t[667] ^ x[117];
  assign t[605] = t[668] ^ x[118];
  assign t[606] = t[669] ^ x[119];
  assign t[607] = t[670] ^ x[120];
  assign t[608] = t[671] ^ x[121];
  assign t[609] = t[672] ^ x[122];
  assign t[60] = ~(t[94] | t[95]);
  assign t[610] = t[673] ^ x[123];
  assign t[611] = t[674] ^ x[124];
  assign t[612] = t[675] ^ x[125];
  assign t[613] = t[676] ^ x[141];
  assign t[614] = t[677] ^ x[157];
  assign t[615] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[616] = (x[0]);
  assign t[617] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[618] = (x[11]);
  assign t[619] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = ~(t[418] | t[96]);
  assign t[620] = (x[14]);
  assign t[621] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[622] = (x[17]);
  assign t[623] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[624] = (x[20]);
  assign t[625] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[626] = (x[24]);
  assign t[627] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[628] = (x[30]);
  assign t[629] = (x[25]);
  assign t[62] = ~(t[97] ^ t[98]);
  assign t[630] = (x[26]);
  assign t[631] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[632] = (x[38]);
  assign t[633] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[634] = (x[46]);
  assign t[635] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[636] = (x[52]);
  assign t[637] = (x[31]);
  assign t[638] = (x[32]);
  assign t[639] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[63] = ~(t[99] | t[100]);
  assign t[640] = (x[60]);
  assign t[641] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[642] = (x[68]);
  assign t[643] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[644] = (x[74]);
  assign t[645] = (x[23]);
  assign t[646] = (x[39]);
  assign t[647] = (x[40]);
  assign t[648] = (x[47]);
  assign t[649] = (x[48]);
  assign t[64] = ~(t[419] | t[101]);
  assign t[650] = (x[53]);
  assign t[651] = (x[54]);
  assign t[652] = (x[88] & ~x[89] & ~x[90] & ~x[91]) | (~x[88] & x[89] & ~x[90] & ~x[91]) | (~x[88] & ~x[89] & x[90] & ~x[91]) | (~x[88] & ~x[89] & ~x[90] & x[91]) | (x[88] & x[89] & x[90] & ~x[91]) | (x[88] & x[89] & ~x[90] & x[91]) | (x[88] & ~x[89] & x[90] & x[91]) | (~x[88] & x[89] & x[90] & x[91]);
  assign t[653] = (x[89]);
  assign t[654] = (x[29]);
  assign t[655] = (x[61]);
  assign t[656] = (x[62]);
  assign t[657] = (x[69]);
  assign t[658] = (x[70]);
  assign t[659] = (x[75]);
  assign t[65] = ~(t[102] | t[103]);
  assign t[660] = (x[76]);
  assign t[661] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[662] = (x[106]);
  assign t[663] = (x[37]);
  assign t[664] = (x[45]);
  assign t[665] = (x[51]);
  assign t[666] = (x[90]);
  assign t[667] = (x[91]);
  assign t[668] = (x[59]);
  assign t[669] = (x[67]);
  assign t[66] = ~(t[104] ^ t[105]);
  assign t[670] = (x[73]);
  assign t[671] = (x[107]);
  assign t[672] = (x[108]);
  assign t[673] = (x[88]);
  assign t[674] = (x[105]);
  assign t[675] = (x[1]);
  assign t[676] = (x[2]);
  assign t[677] = (x[3]);
  assign t[67] = ~(t[420]);
  assign t[68] = ~(t[421]);
  assign t[69] = ~(t[106] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[422] | t[110]);
  assign t[72] = t[111] ? x[66] : x[65];
  assign t[73] = ~(t[112] & t[113]);
  assign t[74] = ~(t[114] | t[115]);
  assign t[75] = ~(t[423] | t[116]);
  assign t[76] = ~(t[117] ^ t[118]);
  assign t[77] = ~(t[119] | t[120]);
  assign t[78] = ~(t[424] | t[121]);
  assign t[79] = ~(t[122] | t[123]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[124] ^ t[125]);
  assign t[81] = ~(t[126]);
  assign t[82] = t[409] ? t[128] : t[127];
  assign t[83] = ~(t[129] | t[130]);
  assign t[84] = ~(t[131] | t[132]);
  assign t[85] = t[409] ? t[134] : t[133];
  assign t[86] = ~(t[425]);
  assign t[87] = ~(t[415] | t[416]);
  assign t[88] = ~(t[426]);
  assign t[89] = ~(t[427]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[135] | t[136]);
  assign t[91] = ~(t[49]);
  assign t[92] = ~(t[129] | t[137]);
  assign t[93] = ~(t[138] | t[139]);
  assign t[94] = ~(t[428]);
  assign t[95] = ~(t[429]);
  assign t[96] = ~(t[140] | t[141]);
  assign t[97] = t[91] ? x[85] : x[84];
  assign t[98] = ~(t[142] & t[143]);
  assign t[99] = ~(t[430]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[211] & ~t[280] & ~t[359]) | (~t[0] & t[211] & ~t[280] & ~t[359]) | (~t[0] & ~t[211] & t[280] & ~t[359]) | (~t[0] & ~t[211] & ~t[280] & t[359]) | (t[0] & t[211] & t[280] & ~t[359]) | (t[0] & t[211] & ~t[280] & t[359]) | (t[0] & ~t[211] & t[280] & t[359]) | (~t[0] & t[211] & t[280] & t[359]);
endmodule

module R2ind171(x, y);
 input [124:0] x;
 output y;

 wire [364:0] t;
  assign t[0] = t[1] ? t[2] : t[110];
  assign t[100] = ~(t[108] | t[98]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[148]);
  assign t[103] = ~(t[149]);
  assign t[104] = ~(t[150]);
  assign t[105] = ~(t[151]);
  assign t[106] = ~(t[152]);
  assign t[107] = ~(t[109] | t[105]);
  assign t[108] = ~(t[153]);
  assign t[109] = ~(t[154]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[155]);
  assign t[111] = (t[156]);
  assign t[112] = (t[157]);
  assign t[113] = (t[158]);
  assign t[114] = (t[159]);
  assign t[115] = (t[160]);
  assign t[116] = (t[161]);
  assign t[117] = (t[162]);
  assign t[118] = (t[163]);
  assign t[119] = (t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = t[200] ^ x[5];
  assign t[156] = t[201] ^ x[13];
  assign t[157] = t[202] ^ x[16];
  assign t[158] = t[203] ^ x[19];
  assign t[159] = t[204] ^ x[22];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[205] ^ x[28];
  assign t[161] = t[206] ^ x[36];
  assign t[162] = t[207] ^ x[39];
  assign t[163] = t[208] ^ x[40];
  assign t[164] = t[209] ^ x[46];
  assign t[165] = t[210] ^ x[52];
  assign t[166] = t[211] ^ x[60];
  assign t[167] = t[212] ^ x[63];
  assign t[168] = t[213] ^ x[64];
  assign t[169] = t[214] ^ x[70];
  assign t[16] = ~(t[111] & t[112]);
  assign t[170] = t[215] ^ x[76];
  assign t[171] = t[216] ^ x[84];
  assign t[172] = t[217] ^ x[87];
  assign t[173] = t[218] ^ x[88];
  assign t[174] = t[219] ^ x[89];
  assign t[175] = t[220] ^ x[90];
  assign t[176] = t[221] ^ x[91];
  assign t[177] = t[222] ^ x[97];
  assign t[178] = t[223] ^ x[98];
  assign t[179] = t[224] ^ x[99];
  assign t[17] = ~(t[113] & t[114]);
  assign t[180] = t[225] ^ x[100];
  assign t[181] = t[226] ^ x[101];
  assign t[182] = t[227] ^ x[102];
  assign t[183] = t[228] ^ x[103];
  assign t[184] = t[229] ^ x[104];
  assign t[185] = t[230] ^ x[105];
  assign t[186] = t[231] ^ x[106];
  assign t[187] = t[232] ^ x[112];
  assign t[188] = t[233] ^ x[113];
  assign t[189] = t[234] ^ x[114];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[115];
  assign t[191] = t[236] ^ x[116];
  assign t[192] = t[237] ^ x[117];
  assign t[193] = t[238] ^ x[118];
  assign t[194] = t[239] ^ x[119];
  assign t[195] = t[240] ^ x[120];
  assign t[196] = t[241] ^ x[121];
  assign t[197] = t[242] ^ x[122];
  assign t[198] = t[243] ^ x[123];
  assign t[199] = t[244] ^ x[124];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[245] & t[246]);
  assign t[201] = (~t[247] & t[248]);
  assign t[202] = (~t[249] & t[250]);
  assign t[203] = (~t[251] & t[252]);
  assign t[204] = (~t[253] & t[254]);
  assign t[205] = (~t[255] & t[256]);
  assign t[206] = (~t[257] & t[258]);
  assign t[207] = (~t[255] & t[259]);
  assign t[208] = (~t[255] & t[260]);
  assign t[209] = (~t[261] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[263] & t[264]);
  assign t[211] = (~t[265] & t[266]);
  assign t[212] = (~t[257] & t[267]);
  assign t[213] = (~t[257] & t[268]);
  assign t[214] = (~t[269] & t[270]);
  assign t[215] = (~t[271] & t[272]);
  assign t[216] = (~t[273] & t[274]);
  assign t[217] = (~t[255] & t[275]);
  assign t[218] = (~t[261] & t[276]);
  assign t[219] = (~t[261] & t[277]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[263] & t[278]);
  assign t[221] = (~t[263] & t[279]);
  assign t[222] = (~t[280] & t[281]);
  assign t[223] = (~t[265] & t[282]);
  assign t[224] = (~t[265] & t[283]);
  assign t[225] = (~t[257] & t[284]);
  assign t[226] = (~t[269] & t[285]);
  assign t[227] = (~t[269] & t[286]);
  assign t[228] = (~t[271] & t[287]);
  assign t[229] = (~t[271] & t[288]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[273] & t[289]);
  assign t[231] = (~t[273] & t[290]);
  assign t[232] = (~t[291] & t[292]);
  assign t[233] = (~t[261] & t[293]);
  assign t[234] = (~t[263] & t[294]);
  assign t[235] = (~t[280] & t[295]);
  assign t[236] = (~t[280] & t[296]);
  assign t[237] = (~t[265] & t[297]);
  assign t[238] = (~t[269] & t[298]);
  assign t[239] = (~t[271] & t[299]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[273] & t[300]);
  assign t[241] = (~t[291] & t[301]);
  assign t[242] = (~t[291] & t[302]);
  assign t[243] = (~t[280] & t[303]);
  assign t[244] = (~t[291] & t[304]);
  assign t[245] = t[305] ^ x[4];
  assign t[246] = t[306] ^ x[5];
  assign t[247] = t[307] ^ x[12];
  assign t[248] = t[308] ^ x[13];
  assign t[249] = t[309] ^ x[15];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[310] ^ x[16];
  assign t[251] = t[311] ^ x[18];
  assign t[252] = t[312] ^ x[19];
  assign t[253] = t[313] ^ x[21];
  assign t[254] = t[314] ^ x[22];
  assign t[255] = t[315] ^ x[27];
  assign t[256] = t[316] ^ x[28];
  assign t[257] = t[317] ^ x[35];
  assign t[258] = t[318] ^ x[36];
  assign t[259] = t[319] ^ x[39];
  assign t[25] = ~(t[113]);
  assign t[260] = t[320] ^ x[40];
  assign t[261] = t[321] ^ x[45];
  assign t[262] = t[322] ^ x[46];
  assign t[263] = t[323] ^ x[51];
  assign t[264] = t[324] ^ x[52];
  assign t[265] = t[325] ^ x[59];
  assign t[266] = t[326] ^ x[60];
  assign t[267] = t[327] ^ x[63];
  assign t[268] = t[328] ^ x[64];
  assign t[269] = t[329] ^ x[69];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[70];
  assign t[271] = t[331] ^ x[75];
  assign t[272] = t[332] ^ x[76];
  assign t[273] = t[333] ^ x[83];
  assign t[274] = t[334] ^ x[84];
  assign t[275] = t[335] ^ x[87];
  assign t[276] = t[336] ^ x[88];
  assign t[277] = t[337] ^ x[89];
  assign t[278] = t[338] ^ x[90];
  assign t[279] = t[339] ^ x[91];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[96];
  assign t[281] = t[341] ^ x[97];
  assign t[282] = t[342] ^ x[98];
  assign t[283] = t[343] ^ x[99];
  assign t[284] = t[344] ^ x[100];
  assign t[285] = t[345] ^ x[101];
  assign t[286] = t[346] ^ x[102];
  assign t[287] = t[347] ^ x[103];
  assign t[288] = t[348] ^ x[104];
  assign t[289] = t[349] ^ x[105];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[106];
  assign t[291] = t[351] ^ x[111];
  assign t[292] = t[352] ^ x[112];
  assign t[293] = t[353] ^ x[113];
  assign t[294] = t[354] ^ x[114];
  assign t[295] = t[355] ^ x[115];
  assign t[296] = t[356] ^ x[116];
  assign t[297] = t[357] ^ x[117];
  assign t[298] = t[358] ^ x[118];
  assign t[299] = t[359] ^ x[119];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[120];
  assign t[301] = t[361] ^ x[121];
  assign t[302] = t[362] ^ x[122];
  assign t[303] = t[363] ^ x[123];
  assign t[304] = t[364] ^ x[124];
  assign t[305] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[306] = (x[3]);
  assign t[307] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[308] = (x[11]);
  assign t[309] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = (x[14]);
  assign t[311] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[312] = (x[17]);
  assign t[313] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[314] = (x[20]);
  assign t[315] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[316] = (x[24]);
  assign t[317] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[318] = (x[32]);
  assign t[319] = (x[26]);
  assign t[31] = t[48] | t[115];
  assign t[320] = (x[23]);
  assign t[321] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[322] = (x[42]);
  assign t[323] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[324] = (x[48]);
  assign t[325] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[326] = (x[56]);
  assign t[327] = (x[34]);
  assign t[328] = (x[31]);
  assign t[329] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[32] = t[49] ? x[30] : x[29];
  assign t[330] = (x[66]);
  assign t[331] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[332] = (x[72]);
  assign t[333] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[334] = (x[80]);
  assign t[335] = (x[25]);
  assign t[336] = (x[44]);
  assign t[337] = (x[41]);
  assign t[338] = (x[50]);
  assign t[339] = (x[47]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[92] & ~x[93] & ~x[94] & ~x[95]) | (~x[92] & x[93] & ~x[94] & ~x[95]) | (~x[92] & ~x[93] & x[94] & ~x[95]) | (~x[92] & ~x[93] & ~x[94] & x[95]) | (x[92] & x[93] & x[94] & ~x[95]) | (x[92] & x[93] & ~x[94] & x[95]) | (x[92] & ~x[93] & x[94] & x[95]) | (~x[92] & x[93] & x[94] & x[95]);
  assign t[341] = (x[93]);
  assign t[342] = (x[58]);
  assign t[343] = (x[55]);
  assign t[344] = (x[33]);
  assign t[345] = (x[68]);
  assign t[346] = (x[65]);
  assign t[347] = (x[74]);
  assign t[348] = (x[71]);
  assign t[349] = (x[82]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[79]);
  assign t[351] = (x[107] & ~x[108] & ~x[109] & ~x[110]) | (~x[107] & x[108] & ~x[109] & ~x[110]) | (~x[107] & ~x[108] & x[109] & ~x[110]) | (~x[107] & ~x[108] & ~x[109] & x[110]) | (x[107] & x[108] & x[109] & ~x[110]) | (x[107] & x[108] & ~x[109] & x[110]) | (x[107] & ~x[108] & x[109] & x[110]) | (~x[107] & x[108] & x[109] & x[110]);
  assign t[352] = (x[108]);
  assign t[353] = (x[43]);
  assign t[354] = (x[49]);
  assign t[355] = (x[95]);
  assign t[356] = (x[92]);
  assign t[357] = (x[57]);
  assign t[358] = (x[67]);
  assign t[359] = (x[73]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[81]);
  assign t[361] = (x[110]);
  assign t[362] = (x[107]);
  assign t[363] = (x[94]);
  assign t[364] = (x[109]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[37] = t[58] ^ t[44];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = t[61] | t[116];
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ? x[38] : x[37];
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[117]);
  assign t[47] = ~(t[118]);
  assign t[48] = ~(t[72] | t[46]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[73] & t[74]);
  assign t[51] = t[75] | t[119];
  assign t[52] = ~(t[76] & t[77]);
  assign t[53] = t[78] | t[120];
  assign t[54] = t[49] ? x[54] : x[53];
  assign t[55] = ~(t[79] & t[80]);
  assign t[56] = ~(t[81] & t[82]);
  assign t[57] = t[83] | t[121];
  assign t[58] = t[62] ? x[62] : x[61];
  assign t[59] = ~(t[122]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[123]);
  assign t[61] = ~(t[84] | t[59]);
  assign t[62] = ~(t[25]);
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = t[87] | t[124];
  assign t[65] = ~(t[88] & t[89]);
  assign t[66] = t[90] | t[125];
  assign t[67] = t[62] ? x[78] : x[77];
  assign t[68] = ~(t[91] & t[92]);
  assign t[69] = t[93] | t[126];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[62] ? x[86] : x[85];
  assign t[71] = ~(t[94] & t[95]);
  assign t[72] = ~(t[127]);
  assign t[73] = ~(t[128]);
  assign t[74] = ~(t[129]);
  assign t[75] = ~(t[96] | t[73]);
  assign t[76] = ~(t[130]);
  assign t[77] = ~(t[131]);
  assign t[78] = ~(t[97] | t[76]);
  assign t[79] = ~(t[98] & t[99]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = t[100] | t[132];
  assign t[81] = ~(t[133]);
  assign t[82] = ~(t[134]);
  assign t[83] = ~(t[101] | t[81]);
  assign t[84] = ~(t[135]);
  assign t[85] = ~(t[136]);
  assign t[86] = ~(t[137]);
  assign t[87] = ~(t[102] | t[85]);
  assign t[88] = ~(t[138]);
  assign t[89] = ~(t[139]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[103] | t[88]);
  assign t[91] = ~(t[140]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[104] | t[91]);
  assign t[94] = ~(t[105] & t[106]);
  assign t[95] = t[107] | t[142];
  assign t[96] = ~(t[143]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[145]);
  assign t[99] = ~(t[146]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [124:0] x;
 output y;

 wire [374:0] t;
  assign t[0] = t[1] ? t[2] : t[120];
  assign t[100] = ~(t[141] & t[140]);
  assign t[101] = ~(t[154]);
  assign t[102] = ~(t[155]);
  assign t[103] = ~(t[156]);
  assign t[104] = ~(t[116] & t[117]);
  assign t[105] = ~(t[144] & t[143]);
  assign t[106] = ~(t[157]);
  assign t[107] = ~(t[147] & t[146]);
  assign t[108] = ~(t[158]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[159]);
  assign t[111] = ~(t[151] & t[150]);
  assign t[112] = ~(t[160]);
  assign t[113] = ~(t[161]);
  assign t[114] = ~(t[162]);
  assign t[115] = ~(t[118] & t[119]);
  assign t[116] = ~(t[156] & t[155]);
  assign t[117] = ~(t[163]);
  assign t[118] = ~(t[162] & t[161]);
  assign t[119] = ~(t[164]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[165]);
  assign t[121] = (t[166]);
  assign t[122] = (t[167]);
  assign t[123] = (t[168]);
  assign t[124] = (t[169]);
  assign t[125] = (t[170]);
  assign t[126] = (t[171]);
  assign t[127] = (t[172]);
  assign t[128] = (t[173]);
  assign t[129] = (t[174]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[175]);
  assign t[131] = (t[176]);
  assign t[132] = (t[177]);
  assign t[133] = (t[178]);
  assign t[134] = (t[179]);
  assign t[135] = (t[180]);
  assign t[136] = (t[181]);
  assign t[137] = (t[182]);
  assign t[138] = (t[183]);
  assign t[139] = (t[184]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[185]);
  assign t[141] = (t[186]);
  assign t[142] = (t[187]);
  assign t[143] = (t[188]);
  assign t[144] = (t[189]);
  assign t[145] = (t[190]);
  assign t[146] = (t[191]);
  assign t[147] = (t[192]);
  assign t[148] = (t[193]);
  assign t[149] = (t[194]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[195]);
  assign t[151] = (t[196]);
  assign t[152] = (t[197]);
  assign t[153] = (t[198]);
  assign t[154] = (t[199]);
  assign t[155] = (t[200]);
  assign t[156] = (t[201]);
  assign t[157] = (t[202]);
  assign t[158] = (t[203]);
  assign t[159] = (t[204]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (t[205]);
  assign t[161] = (t[206]);
  assign t[162] = (t[207]);
  assign t[163] = (t[208]);
  assign t[164] = (t[209]);
  assign t[165] = t[210] ^ x[5];
  assign t[166] = t[211] ^ x[13];
  assign t[167] = t[212] ^ x[16];
  assign t[168] = t[213] ^ x[19];
  assign t[169] = t[214] ^ x[22];
  assign t[16] = ~(t[121] & t[122]);
  assign t[170] = t[215] ^ x[28];
  assign t[171] = t[216] ^ x[36];
  assign t[172] = t[217] ^ x[39];
  assign t[173] = t[218] ^ x[40];
  assign t[174] = t[219] ^ x[46];
  assign t[175] = t[220] ^ x[52];
  assign t[176] = t[221] ^ x[60];
  assign t[177] = t[222] ^ x[63];
  assign t[178] = t[223] ^ x[64];
  assign t[179] = t[224] ^ x[70];
  assign t[17] = ~(t[123] & t[124]);
  assign t[180] = t[225] ^ x[76];
  assign t[181] = t[226] ^ x[84];
  assign t[182] = t[227] ^ x[87];
  assign t[183] = t[228] ^ x[88];
  assign t[184] = t[229] ^ x[89];
  assign t[185] = t[230] ^ x[90];
  assign t[186] = t[231] ^ x[91];
  assign t[187] = t[232] ^ x[97];
  assign t[188] = t[233] ^ x[98];
  assign t[189] = t[234] ^ x[99];
  assign t[18] = ~(t[25]);
  assign t[190] = t[235] ^ x[100];
  assign t[191] = t[236] ^ x[101];
  assign t[192] = t[237] ^ x[102];
  assign t[193] = t[238] ^ x[103];
  assign t[194] = t[239] ^ x[104];
  assign t[195] = t[240] ^ x[105];
  assign t[196] = t[241] ^ x[106];
  assign t[197] = t[242] ^ x[112];
  assign t[198] = t[243] ^ x[113];
  assign t[199] = t[244] ^ x[114];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[245] ^ x[115];
  assign t[201] = t[246] ^ x[116];
  assign t[202] = t[247] ^ x[117];
  assign t[203] = t[248] ^ x[118];
  assign t[204] = t[249] ^ x[119];
  assign t[205] = t[250] ^ x[120];
  assign t[206] = t[251] ^ x[121];
  assign t[207] = t[252] ^ x[122];
  assign t[208] = t[253] ^ x[123];
  assign t[209] = t[254] ^ x[124];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[255] & t[256]);
  assign t[211] = (~t[257] & t[258]);
  assign t[212] = (~t[259] & t[260]);
  assign t[213] = (~t[261] & t[262]);
  assign t[214] = (~t[263] & t[264]);
  assign t[215] = (~t[265] & t[266]);
  assign t[216] = (~t[267] & t[268]);
  assign t[217] = (~t[265] & t[269]);
  assign t[218] = (~t[265] & t[270]);
  assign t[219] = (~t[271] & t[272]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[273] & t[274]);
  assign t[221] = (~t[275] & t[276]);
  assign t[222] = (~t[267] & t[277]);
  assign t[223] = (~t[267] & t[278]);
  assign t[224] = (~t[279] & t[280]);
  assign t[225] = (~t[281] & t[282]);
  assign t[226] = (~t[283] & t[284]);
  assign t[227] = (~t[265] & t[285]);
  assign t[228] = (~t[271] & t[286]);
  assign t[229] = (~t[271] & t[287]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[273] & t[288]);
  assign t[231] = (~t[273] & t[289]);
  assign t[232] = (~t[290] & t[291]);
  assign t[233] = (~t[275] & t[292]);
  assign t[234] = (~t[275] & t[293]);
  assign t[235] = (~t[267] & t[294]);
  assign t[236] = (~t[279] & t[295]);
  assign t[237] = (~t[279] & t[296]);
  assign t[238] = (~t[281] & t[297]);
  assign t[239] = (~t[281] & t[298]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (~t[283] & t[299]);
  assign t[241] = (~t[283] & t[300]);
  assign t[242] = (~t[301] & t[302]);
  assign t[243] = (~t[271] & t[303]);
  assign t[244] = (~t[273] & t[304]);
  assign t[245] = (~t[290] & t[305]);
  assign t[246] = (~t[290] & t[306]);
  assign t[247] = (~t[275] & t[307]);
  assign t[248] = (~t[279] & t[308]);
  assign t[249] = (~t[281] & t[309]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = (~t[283] & t[310]);
  assign t[251] = (~t[301] & t[311]);
  assign t[252] = (~t[301] & t[312]);
  assign t[253] = (~t[290] & t[313]);
  assign t[254] = (~t[301] & t[314]);
  assign t[255] = t[315] ^ x[4];
  assign t[256] = t[316] ^ x[5];
  assign t[257] = t[317] ^ x[12];
  assign t[258] = t[318] ^ x[13];
  assign t[259] = t[319] ^ x[15];
  assign t[25] = ~(t[123]);
  assign t[260] = t[320] ^ x[16];
  assign t[261] = t[321] ^ x[18];
  assign t[262] = t[322] ^ x[19];
  assign t[263] = t[323] ^ x[21];
  assign t[264] = t[324] ^ x[22];
  assign t[265] = t[325] ^ x[27];
  assign t[266] = t[326] ^ x[28];
  assign t[267] = t[327] ^ x[35];
  assign t[268] = t[328] ^ x[36];
  assign t[269] = t[329] ^ x[39];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[330] ^ x[40];
  assign t[271] = t[331] ^ x[45];
  assign t[272] = t[332] ^ x[46];
  assign t[273] = t[333] ^ x[51];
  assign t[274] = t[334] ^ x[52];
  assign t[275] = t[335] ^ x[59];
  assign t[276] = t[336] ^ x[60];
  assign t[277] = t[337] ^ x[63];
  assign t[278] = t[338] ^ x[64];
  assign t[279] = t[339] ^ x[69];
  assign t[27] = t[40] ^ t[41];
  assign t[280] = t[340] ^ x[70];
  assign t[281] = t[341] ^ x[75];
  assign t[282] = t[342] ^ x[76];
  assign t[283] = t[343] ^ x[83];
  assign t[284] = t[344] ^ x[84];
  assign t[285] = t[345] ^ x[87];
  assign t[286] = t[346] ^ x[88];
  assign t[287] = t[347] ^ x[89];
  assign t[288] = t[348] ^ x[90];
  assign t[289] = t[349] ^ x[91];
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = t[350] ^ x[96];
  assign t[291] = t[351] ^ x[97];
  assign t[292] = t[352] ^ x[98];
  assign t[293] = t[353] ^ x[99];
  assign t[294] = t[354] ^ x[100];
  assign t[295] = t[355] ^ x[101];
  assign t[296] = t[356] ^ x[102];
  assign t[297] = t[357] ^ x[103];
  assign t[298] = t[358] ^ x[104];
  assign t[299] = t[359] ^ x[105];
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[360] ^ x[106];
  assign t[301] = t[361] ^ x[111];
  assign t[302] = t[362] ^ x[112];
  assign t[303] = t[363] ^ x[113];
  assign t[304] = t[364] ^ x[114];
  assign t[305] = t[365] ^ x[115];
  assign t[306] = t[366] ^ x[116];
  assign t[307] = t[367] ^ x[117];
  assign t[308] = t[368] ^ x[118];
  assign t[309] = t[369] ^ x[119];
  assign t[30] = ~(t[46] & t[47]);
  assign t[310] = t[370] ^ x[120];
  assign t[311] = t[371] ^ x[121];
  assign t[312] = t[372] ^ x[122];
  assign t[313] = t[373] ^ x[123];
  assign t[314] = t[374] ^ x[124];
  assign t[315] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[316] = (x[2]);
  assign t[317] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[318] = (x[11]);
  assign t[319] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = ~(t[48] & t[125]);
  assign t[320] = (x[14]);
  assign t[321] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[322] = (x[17]);
  assign t[323] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[324] = (x[20]);
  assign t[325] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[326] = (x[24]);
  assign t[327] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[328] = (x[32]);
  assign t[329] = (x[26]);
  assign t[32] = t[49] ? x[30] : x[29];
  assign t[330] = (x[23]);
  assign t[331] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[332] = (x[42]);
  assign t[333] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[334] = (x[48]);
  assign t[335] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[336] = (x[56]);
  assign t[337] = (x[34]);
  assign t[338] = (x[31]);
  assign t[339] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[33] = ~(t[50] & t[51]);
  assign t[340] = (x[66]);
  assign t[341] = (x[71] & ~x[72] & ~x[73] & ~x[74]) | (~x[71] & x[72] & ~x[73] & ~x[74]) | (~x[71] & ~x[72] & x[73] & ~x[74]) | (~x[71] & ~x[72] & ~x[73] & x[74]) | (x[71] & x[72] & x[73] & ~x[74]) | (x[71] & x[72] & ~x[73] & x[74]) | (x[71] & ~x[72] & x[73] & x[74]) | (~x[71] & x[72] & x[73] & x[74]);
  assign t[342] = (x[72]);
  assign t[343] = (x[79] & ~x[80] & ~x[81] & ~x[82]) | (~x[79] & x[80] & ~x[81] & ~x[82]) | (~x[79] & ~x[80] & x[81] & ~x[82]) | (~x[79] & ~x[80] & ~x[81] & x[82]) | (x[79] & x[80] & x[81] & ~x[82]) | (x[79] & x[80] & ~x[81] & x[82]) | (x[79] & ~x[80] & x[81] & x[82]) | (~x[79] & x[80] & x[81] & x[82]);
  assign t[344] = (x[80]);
  assign t[345] = (x[25]);
  assign t[346] = (x[44]);
  assign t[347] = (x[41]);
  assign t[348] = (x[50]);
  assign t[349] = (x[47]);
  assign t[34] = ~(t[52] & t[53]);
  assign t[350] = (x[92] & ~x[93] & ~x[94] & ~x[95]) | (~x[92] & x[93] & ~x[94] & ~x[95]) | (~x[92] & ~x[93] & x[94] & ~x[95]) | (~x[92] & ~x[93] & ~x[94] & x[95]) | (x[92] & x[93] & x[94] & ~x[95]) | (x[92] & x[93] & ~x[94] & x[95]) | (x[92] & ~x[93] & x[94] & x[95]) | (~x[92] & x[93] & x[94] & x[95]);
  assign t[351] = (x[93]);
  assign t[352] = (x[58]);
  assign t[353] = (x[55]);
  assign t[354] = (x[33]);
  assign t[355] = (x[68]);
  assign t[356] = (x[65]);
  assign t[357] = (x[74]);
  assign t[358] = (x[71]);
  assign t[359] = (x[82]);
  assign t[35] = t[54] ^ t[55];
  assign t[360] = (x[79]);
  assign t[361] = (x[107] & ~x[108] & ~x[109] & ~x[110]) | (~x[107] & x[108] & ~x[109] & ~x[110]) | (~x[107] & ~x[108] & x[109] & ~x[110]) | (~x[107] & ~x[108] & ~x[109] & x[110]) | (x[107] & x[108] & x[109] & ~x[110]) | (x[107] & x[108] & ~x[109] & x[110]) | (x[107] & ~x[108] & x[109] & x[110]) | (~x[107] & x[108] & x[109] & x[110]);
  assign t[362] = (x[108]);
  assign t[363] = (x[43]);
  assign t[364] = (x[49]);
  assign t[365] = (x[95]);
  assign t[366] = (x[92]);
  assign t[367] = (x[57]);
  assign t[368] = (x[67]);
  assign t[369] = (x[73]);
  assign t[36] = ~(t[56] & t[57]);
  assign t[370] = (x[81]);
  assign t[371] = (x[110]);
  assign t[372] = (x[107]);
  assign t[373] = (x[94]);
  assign t[374] = (x[109]);
  assign t[37] = t[58] ^ t[44];
  assign t[38] = ~(t[59] & t[60]);
  assign t[39] = ~(t[61] & t[126]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ? x[38] : x[37];
  assign t[41] = ~(t[63] & t[64]);
  assign t[42] = ~(t[65] & t[66]);
  assign t[43] = t[67] ^ t[42];
  assign t[44] = ~(t[68] & t[69]);
  assign t[45] = t[70] ^ t[71];
  assign t[46] = ~(t[127]);
  assign t[47] = ~(t[128]);
  assign t[48] = ~(t[72] & t[73]);
  assign t[49] = ~(t[25]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[74] & t[75]);
  assign t[51] = ~(t[76] & t[129]);
  assign t[52] = ~(t[77] & t[78]);
  assign t[53] = ~(t[79] & t[130]);
  assign t[54] = t[49] ? x[54] : x[53];
  assign t[55] = ~(t[80] & t[81]);
  assign t[56] = ~(t[82] & t[83]);
  assign t[57] = ~(t[84] & t[131]);
  assign t[58] = t[18] ? x[62] : x[61];
  assign t[59] = ~(t[132]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[133]);
  assign t[61] = ~(t[85] & t[86]);
  assign t[62] = ~(t[25]);
  assign t[63] = ~(t[87] & t[88]);
  assign t[64] = ~(t[89] & t[134]);
  assign t[65] = ~(t[90] & t[91]);
  assign t[66] = ~(t[92] & t[135]);
  assign t[67] = t[62] ? x[78] : x[77];
  assign t[68] = ~(t[93] & t[94]);
  assign t[69] = ~(t[95] & t[136]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[62] ? x[86] : x[85];
  assign t[71] = ~(t[96] & t[97]);
  assign t[72] = ~(t[128] & t[127]);
  assign t[73] = ~(t[137]);
  assign t[74] = ~(t[138]);
  assign t[75] = ~(t[139]);
  assign t[76] = ~(t[98] & t[99]);
  assign t[77] = ~(t[140]);
  assign t[78] = ~(t[141]);
  assign t[79] = ~(t[100] & t[101]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[102] & t[103]);
  assign t[81] = ~(t[104] & t[142]);
  assign t[82] = ~(t[143]);
  assign t[83] = ~(t[144]);
  assign t[84] = ~(t[105] & t[106]);
  assign t[85] = ~(t[133] & t[132]);
  assign t[86] = ~(t[145]);
  assign t[87] = ~(t[146]);
  assign t[88] = ~(t[147]);
  assign t[89] = ~(t[107] & t[108]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[148]);
  assign t[91] = ~(t[149]);
  assign t[92] = ~(t[109] & t[110]);
  assign t[93] = ~(t[150]);
  assign t[94] = ~(t[151]);
  assign t[95] = ~(t[111] & t[112]);
  assign t[96] = ~(t[113] & t[114]);
  assign t[97] = ~(t[115] & t[152]);
  assign t[98] = ~(t[139] & t[138]);
  assign t[99] = ~(t[153]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [114:0] x;
 output y;

 wire [304:0] t;
  assign t[0] = t[1] ? t[2] : t[100];
  assign t[100] = (t[135]);
  assign t[101] = (t[136]);
  assign t[102] = (t[137]);
  assign t[103] = (t[138]);
  assign t[104] = (t[139]);
  assign t[105] = (t[140]);
  assign t[106] = (t[141]);
  assign t[107] = (t[142]);
  assign t[108] = (t[143]);
  assign t[109] = (t[144]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[145]);
  assign t[111] = (t[146]);
  assign t[112] = (t[147]);
  assign t[113] = (t[148]);
  assign t[114] = (t[149]);
  assign t[115] = (t[150]);
  assign t[116] = (t[151]);
  assign t[117] = (t[152]);
  assign t[118] = (t[153]);
  assign t[119] = (t[154]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[155]);
  assign t[121] = (t[156]);
  assign t[122] = (t[157]);
  assign t[123] = (t[158]);
  assign t[124] = (t[159]);
  assign t[125] = (t[160]);
  assign t[126] = (t[161]);
  assign t[127] = (t[162]);
  assign t[128] = (t[163]);
  assign t[129] = (t[164]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[165]);
  assign t[131] = (t[166]);
  assign t[132] = (t[167]);
  assign t[133] = (t[168]);
  assign t[134] = (t[169]);
  assign t[135] = t[170] ^ x[5];
  assign t[136] = t[171] ^ x[13];
  assign t[137] = t[172] ^ x[16];
  assign t[138] = t[173] ^ x[19];
  assign t[139] = t[174] ^ x[22];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[175] ^ x[28];
  assign t[141] = t[176] ^ x[29];
  assign t[142] = t[177] ^ x[37];
  assign t[143] = t[178] ^ x[38];
  assign t[144] = t[179] ^ x[41];
  assign t[145] = t[180] ^ x[47];
  assign t[146] = t[181] ^ x[48];
  assign t[147] = t[182] ^ x[54];
  assign t[148] = t[183] ^ x[55];
  assign t[149] = t[184] ^ x[63];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[185] ^ x[64];
  assign t[151] = t[186] ^ x[67];
  assign t[152] = t[187] ^ x[73];
  assign t[153] = t[188] ^ x[74];
  assign t[154] = t[189] ^ x[80];
  assign t[155] = t[190] ^ x[81];
  assign t[156] = t[191] ^ x[89];
  assign t[157] = t[192] ^ x[90];
  assign t[158] = t[193] ^ x[93];
  assign t[159] = t[194] ^ x[94];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[195] ^ x[100];
  assign t[161] = t[196] ^ x[101];
  assign t[162] = t[197] ^ x[102];
  assign t[163] = t[198] ^ x[103];
  assign t[164] = t[199] ^ x[104];
  assign t[165] = t[200] ^ x[110];
  assign t[166] = t[201] ^ x[111];
  assign t[167] = t[202] ^ x[112];
  assign t[168] = t[203] ^ x[113];
  assign t[169] = t[204] ^ x[114];
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (~t[205] & t[206]);
  assign t[171] = (~t[207] & t[208]);
  assign t[172] = (~t[209] & t[210]);
  assign t[173] = (~t[211] & t[212]);
  assign t[174] = (~t[213] & t[214]);
  assign t[175] = (~t[215] & t[216]);
  assign t[176] = (~t[215] & t[217]);
  assign t[177] = (~t[218] & t[219]);
  assign t[178] = (~t[218] & t[220]);
  assign t[179] = (~t[215] & t[221]);
  assign t[17] = ~(t[103] & t[104]);
  assign t[180] = (~t[222] & t[223]);
  assign t[181] = (~t[222] & t[224]);
  assign t[182] = (~t[225] & t[226]);
  assign t[183] = (~t[225] & t[227]);
  assign t[184] = (~t[228] & t[229]);
  assign t[185] = (~t[228] & t[230]);
  assign t[186] = (~t[218] & t[231]);
  assign t[187] = (~t[232] & t[233]);
  assign t[188] = (~t[232] & t[234]);
  assign t[189] = (~t[235] & t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (~t[235] & t[237]);
  assign t[191] = (~t[238] & t[239]);
  assign t[192] = (~t[238] & t[240]);
  assign t[193] = (~t[222] & t[241]);
  assign t[194] = (~t[225] & t[242]);
  assign t[195] = (~t[243] & t[244]);
  assign t[196] = (~t[243] & t[245]);
  assign t[197] = (~t[228] & t[246]);
  assign t[198] = (~t[232] & t[247]);
  assign t[199] = (~t[235] & t[248]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[249] & t[250]);
  assign t[201] = (~t[249] & t[251]);
  assign t[202] = (~t[238] & t[252]);
  assign t[203] = (~t[243] & t[253]);
  assign t[204] = (~t[249] & t[254]);
  assign t[205] = t[255] ^ x[4];
  assign t[206] = t[256] ^ x[5];
  assign t[207] = t[257] ^ x[12];
  assign t[208] = t[258] ^ x[13];
  assign t[209] = t[259] ^ x[15];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[260] ^ x[16];
  assign t[211] = t[261] ^ x[18];
  assign t[212] = t[262] ^ x[19];
  assign t[213] = t[263] ^ x[21];
  assign t[214] = t[264] ^ x[22];
  assign t[215] = t[265] ^ x[27];
  assign t[216] = t[266] ^ x[28];
  assign t[217] = t[267] ^ x[29];
  assign t[218] = t[268] ^ x[36];
  assign t[219] = t[269] ^ x[37];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[270] ^ x[38];
  assign t[221] = t[271] ^ x[41];
  assign t[222] = t[272] ^ x[46];
  assign t[223] = t[273] ^ x[47];
  assign t[224] = t[274] ^ x[48];
  assign t[225] = t[275] ^ x[53];
  assign t[226] = t[276] ^ x[54];
  assign t[227] = t[277] ^ x[55];
  assign t[228] = t[278] ^ x[62];
  assign t[229] = t[279] ^ x[63];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[280] ^ x[64];
  assign t[231] = t[281] ^ x[67];
  assign t[232] = t[282] ^ x[72];
  assign t[233] = t[283] ^ x[73];
  assign t[234] = t[284] ^ x[74];
  assign t[235] = t[285] ^ x[79];
  assign t[236] = t[286] ^ x[80];
  assign t[237] = t[287] ^ x[81];
  assign t[238] = t[288] ^ x[88];
  assign t[239] = t[289] ^ x[89];
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = t[290] ^ x[90];
  assign t[241] = t[291] ^ x[93];
  assign t[242] = t[292] ^ x[94];
  assign t[243] = t[293] ^ x[99];
  assign t[244] = t[294] ^ x[100];
  assign t[245] = t[295] ^ x[101];
  assign t[246] = t[296] ^ x[102];
  assign t[247] = t[297] ^ x[103];
  assign t[248] = t[298] ^ x[104];
  assign t[249] = t[299] ^ x[109];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[300] ^ x[110];
  assign t[251] = t[301] ^ x[111];
  assign t[252] = t[302] ^ x[112];
  assign t[253] = t[303] ^ x[113];
  assign t[254] = t[304] ^ x[114];
  assign t[255] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[256] = (x[1]);
  assign t[257] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[258] = (x[11]);
  assign t[259] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[25] = ~(t[103]);
  assign t[260] = (x[14]);
  assign t[261] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[262] = (x[17]);
  assign t[263] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[264] = (x[20]);
  assign t[265] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[266] = (x[25]);
  assign t[267] = (x[23]);
  assign t[268] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[269] = (x[34]);
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = (x[32]);
  assign t[271] = (x[26]);
  assign t[272] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[273] = (x[44]);
  assign t[274] = (x[42]);
  assign t[275] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[276] = (x[51]);
  assign t[277] = (x[49]);
  assign t[278] = (x[58] & ~x[59] & ~x[60] & ~x[61]) | (~x[58] & x[59] & ~x[60] & ~x[61]) | (~x[58] & ~x[59] & x[60] & ~x[61]) | (~x[58] & ~x[59] & ~x[60] & x[61]) | (x[58] & x[59] & x[60] & ~x[61]) | (x[58] & x[59] & ~x[60] & x[61]) | (x[58] & ~x[59] & x[60] & x[61]) | (~x[58] & x[59] & x[60] & x[61]);
  assign t[279] = (x[60]);
  assign t[27] = t[40] ^ t[41];
  assign t[280] = (x[58]);
  assign t[281] = (x[35]);
  assign t[282] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[283] = (x[70]);
  assign t[284] = (x[68]);
  assign t[285] = (x[75] & ~x[76] & ~x[77] & ~x[78]) | (~x[75] & x[76] & ~x[77] & ~x[78]) | (~x[75] & ~x[76] & x[77] & ~x[78]) | (~x[75] & ~x[76] & ~x[77] & x[78]) | (x[75] & x[76] & x[77] & ~x[78]) | (x[75] & x[76] & ~x[77] & x[78]) | (x[75] & ~x[76] & x[77] & x[78]) | (~x[75] & x[76] & x[77] & x[78]);
  assign t[286] = (x[77]);
  assign t[287] = (x[75]);
  assign t[288] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[289] = (x[86]);
  assign t[28] = x[7] ? t[43] : t[42];
  assign t[290] = (x[84]);
  assign t[291] = (x[45]);
  assign t[292] = (x[52]);
  assign t[293] = (x[95] & ~x[96] & ~x[97] & ~x[98]) | (~x[95] & x[96] & ~x[97] & ~x[98]) | (~x[95] & ~x[96] & x[97] & ~x[98]) | (~x[95] & ~x[96] & ~x[97] & x[98]) | (x[95] & x[96] & x[97] & ~x[98]) | (x[95] & x[96] & ~x[97] & x[98]) | (x[95] & ~x[96] & x[97] & x[98]) | (~x[95] & x[96] & x[97] & x[98]);
  assign t[294] = (x[97]);
  assign t[295] = (x[95]);
  assign t[296] = (x[61]);
  assign t[297] = (x[71]);
  assign t[298] = (x[78]);
  assign t[299] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[29] = x[7] ? t[45] : t[44];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[107]);
  assign t[301] = (x[105]);
  assign t[302] = (x[87]);
  assign t[303] = (x[98]);
  assign t[304] = (x[108]);
  assign t[30] = ~(t[105] & t[46]);
  assign t[31] = ~(t[106] & t[47]);
  assign t[32] = t[48] ? x[31] : x[30];
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[54];
  assign t[36] = ~(t[55] & t[56]);
  assign t[37] = t[57] ^ t[42];
  assign t[38] = ~(t[107] & t[58]);
  assign t[39] = ~(t[108] & t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ? x[40] : x[39];
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = ~(t[63] & t[64]);
  assign t[43] = t[65] ^ t[66];
  assign t[44] = ~(t[67] & t[68]);
  assign t[45] = t[69] ^ t[44];
  assign t[46] = ~(t[109]);
  assign t[47] = ~(t[109] & t[70]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[110] & t[71]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[111] & t[72]);
  assign t[51] = ~(t[112] & t[73]);
  assign t[52] = ~(t[113] & t[74]);
  assign t[53] = t[60] ? x[57] : x[56];
  assign t[54] = ~(t[75] & t[76]);
  assign t[55] = ~(t[114] & t[77]);
  assign t[56] = ~(t[115] & t[78]);
  assign t[57] = t[48] ? x[66] : x[65];
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[116] & t[79]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[25]);
  assign t[61] = ~(t[117] & t[80]);
  assign t[62] = ~(t[118] & t[81]);
  assign t[63] = ~(t[119] & t[82]);
  assign t[64] = ~(t[120] & t[83]);
  assign t[65] = t[60] ? x[83] : x[82];
  assign t[66] = ~(t[84] & t[85]);
  assign t[67] = ~(t[121] & t[86]);
  assign t[68] = ~(t[122] & t[87]);
  assign t[69] = t[60] ? x[92] : x[91];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105]);
  assign t[71] = ~(t[123]);
  assign t[72] = ~(t[123] & t[88]);
  assign t[73] = ~(t[124]);
  assign t[74] = ~(t[124] & t[89]);
  assign t[75] = ~(t[125] & t[90]);
  assign t[76] = ~(t[126] & t[91]);
  assign t[77] = ~(t[127]);
  assign t[78] = ~(t[127] & t[92]);
  assign t[79] = ~(t[107]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[128]);
  assign t[81] = ~(t[128] & t[93]);
  assign t[82] = ~(t[129]);
  assign t[83] = ~(t[129] & t[94]);
  assign t[84] = ~(t[130] & t[95]);
  assign t[85] = ~(t[131] & t[96]);
  assign t[86] = ~(t[132]);
  assign t[87] = ~(t[132] & t[97]);
  assign t[88] = ~(t[110]);
  assign t[89] = ~(t[112]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[133] & t[98]);
  assign t[92] = ~(t[114]);
  assign t[93] = ~(t[117]);
  assign t[94] = ~(t[119]);
  assign t[95] = ~(t[134]);
  assign t[96] = ~(t[134] & t[99]);
  assign t[97] = ~(t[121]);
  assign t[98] = ~(t[125]);
  assign t[99] = ~(t[130]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [124:0] x;
 output y;

 wire [465:0] t;
  assign t[0] = t[1] ? t[2] : t[211];
  assign t[100] = ~(t[234]);
  assign t[101] = ~(t[144] | t[145]);
  assign t[102] = ~(t[146] | t[147]);
  assign t[103] = ~(t[235] | t[148]);
  assign t[104] = t[91] ? x[95] : x[94];
  assign t[105] = ~(t[149] & t[150]);
  assign t[106] = ~(t[236]);
  assign t[107] = ~(t[223] | t[224]);
  assign t[108] = ~(t[237]);
  assign t[109] = ~(t[238]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151] | t[152]);
  assign t[111] = ~(t[49]);
  assign t[112] = ~(t[137] | t[153]);
  assign t[113] = ~(t[154] | t[155]);
  assign t[114] = ~(t[239]);
  assign t[115] = ~(t[240]);
  assign t[116] = ~(t[156] | t[157]);
  assign t[117] = t[111] ? x[102] : x[101];
  assign t[118] = ~(t[158] & t[159]);
  assign t[119] = ~(t[241]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[242]);
  assign t[121] = ~(t[160] | t[161]);
  assign t[122] = ~(t[162] | t[163]);
  assign t[123] = ~(t[243] | t[164]);
  assign t[124] = t[111] ? x[112] : x[111];
  assign t[125] = ~(t[84] & t[149]);
  assign t[126] = ~(t[214]);
  assign t[127] = ~(t[165] & t[166]);
  assign t[128] = ~(x[7] & t[167]);
  assign t[129] = ~(t[81] | t[168]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[142] & t[169]);
  assign t[131] = ~(t[126] | t[170]);
  assign t[132] = ~(t[126] | t[171]);
  assign t[133] = ~(t[172] & t[215]);
  assign t[134] = ~(t[173] & t[166]);
  assign t[135] = ~(t[244]);
  assign t[136] = ~(t[229] | t[230]);
  assign t[137] = ~(t[81] | t[174]);
  assign t[138] = t[175] | t[176];
  assign t[139] = ~(t[177] & t[178]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[245]);
  assign t[141] = ~(t[231] | t[232]);
  assign t[142] = ~(t[179] | t[180]);
  assign t[143] = ~(t[181] | t[182]);
  assign t[144] = ~(t[246]);
  assign t[145] = ~(t[233] | t[234]);
  assign t[146] = ~(t[247]);
  assign t[147] = ~(t[248]);
  assign t[148] = ~(t[183] | t[184]);
  assign t[149] = ~(t[130] | t[185]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[129] | t[153]);
  assign t[151] = ~(t[249]);
  assign t[152] = ~(t[237] | t[238]);
  assign t[153] = ~(t[81] | t[186]);
  assign t[154] = t[215] & t[187];
  assign t[155] = ~(t[84]);
  assign t[156] = ~(t[250]);
  assign t[157] = ~(t[239] | t[240]);
  assign t[158] = ~(t[179] | t[132]);
  assign t[159] = ~(t[188] | t[176]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = ~(t[251]);
  assign t[161] = ~(t[241] | t[242]);
  assign t[162] = ~(t[252]);
  assign t[163] = ~(t[253]);
  assign t[164] = ~(t[189] | t[190]);
  assign t[165] = ~(x[7] | t[191]);
  assign t[166] = ~(t[215]);
  assign t[167] = ~(t[213] | t[166]);
  assign t[168] = t[212] ? t[133] : t[134];
  assign t[169] = ~(t[126] & t[192]);
  assign t[16] = ~(t[212] & t[213]);
  assign t[170] = t[212] ? t[193] : t[134];
  assign t[171] = t[212] ? t[127] : t[194];
  assign t[172] = x[7] & t[213];
  assign t[173] = ~(x[7] | t[213]);
  assign t[174] = t[212] ? t[194] : t[195];
  assign t[175] = ~(t[84] & t[196]);
  assign t[176] = ~(t[81] | t[197]);
  assign t[177] = ~(t[198] | t[50]);
  assign t[178] = t[126] | t[199];
  assign t[179] = ~(t[126] | t[200]);
  assign t[17] = ~(t[214] & t[215]);
  assign t[180] = ~(t[81] | t[201]);
  assign t[181] = ~(t[81] | t[202]);
  assign t[182] = ~(t[150] & t[178]);
  assign t[183] = ~(t[254]);
  assign t[184] = ~(t[247] | t[248]);
  assign t[185] = ~(t[203] & t[178]);
  assign t[186] = t[212] ? t[193] : t[204];
  assign t[187] = ~(t[126] | t[212]);
  assign t[188] = ~(t[205]);
  assign t[189] = ~(t[255]);
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[252] | t[253]);
  assign t[191] = ~(t[213]);
  assign t[192] = ~(t[194] & t[195]);
  assign t[193] = ~(t[172] & t[166]);
  assign t[194] = ~(x[7] & t[206]);
  assign t[195] = ~(t[215] & t[165]);
  assign t[196] = ~(t[167] & t[207]);
  assign t[197] = t[212] ? t[195] : t[194];
  assign t[198] = ~(t[208]);
  assign t[199] = t[212] ? t[194] : t[127];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[212] ? t[134] : t[193];
  assign t[201] = t[212] ? t[127] : t[128];
  assign t[202] = t[212] ? t[204] : t[193];
  assign t[203] = ~(t[154] & t[209]);
  assign t[204] = ~(t[173] & t[215]);
  assign t[205] = ~(t[50] | t[153]);
  assign t[206] = ~(t[213] | t[215]);
  assign t[207] = t[81] & t[212];
  assign t[208] = ~(t[187] & t[210]);
  assign t[209] = t[173] | t[172];
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = ~(t[195] & t[128]);
  assign t[211] = (t[256]);
  assign t[212] = (t[257]);
  assign t[213] = (t[258]);
  assign t[214] = (t[259]);
  assign t[215] = (t[260]);
  assign t[216] = (t[261]);
  assign t[217] = (t[262]);
  assign t[218] = (t[263]);
  assign t[219] = (t[264]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[265]);
  assign t[221] = (t[266]);
  assign t[222] = (t[267]);
  assign t[223] = (t[268]);
  assign t[224] = (t[269]);
  assign t[225] = (t[270]);
  assign t[226] = (t[271]);
  assign t[227] = (t[272]);
  assign t[228] = (t[273]);
  assign t[229] = (t[274]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[275]);
  assign t[231] = (t[276]);
  assign t[232] = (t[277]);
  assign t[233] = (t[278]);
  assign t[234] = (t[279]);
  assign t[235] = (t[280]);
  assign t[236] = (t[281]);
  assign t[237] = (t[282]);
  assign t[238] = (t[283]);
  assign t[239] = (t[284]);
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = (t[285]);
  assign t[241] = (t[286]);
  assign t[242] = (t[287]);
  assign t[243] = (t[288]);
  assign t[244] = (t[289]);
  assign t[245] = (t[290]);
  assign t[246] = (t[291]);
  assign t[247] = (t[292]);
  assign t[248] = (t[293]);
  assign t[249] = (t[294]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = (t[295]);
  assign t[251] = (t[296]);
  assign t[252] = (t[297]);
  assign t[253] = (t[298]);
  assign t[254] = (t[299]);
  assign t[255] = (t[300]);
  assign t[256] = t[301] ^ x[5];
  assign t[257] = t[302] ^ x[13];
  assign t[258] = t[303] ^ x[16];
  assign t[259] = t[304] ^ x[19];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[305] ^ x[22];
  assign t[261] = t[306] ^ x[28];
  assign t[262] = t[307] ^ x[34];
  assign t[263] = t[308] ^ x[35];
  assign t[264] = t[309] ^ x[36];
  assign t[265] = t[310] ^ x[42];
  assign t[266] = t[311] ^ x[50];
  assign t[267] = t[312] ^ x[56];
  assign t[268] = t[313] ^ x[57];
  assign t[269] = t[314] ^ x[58];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[315] ^ x[64];
  assign t[271] = t[316] ^ x[72];
  assign t[272] = t[317] ^ x[78];
  assign t[273] = t[318] ^ x[79];
  assign t[274] = t[319] ^ x[80];
  assign t[275] = t[320] ^ x[81];
  assign t[276] = t[321] ^ x[82];
  assign t[277] = t[322] ^ x[83];
  assign t[278] = t[323] ^ x[86];
  assign t[279] = t[324] ^ x[87];
  assign t[27] = ~(t[43] ^ t[44]);
  assign t[280] = t[325] ^ x[93];
  assign t[281] = t[326] ^ x[96];
  assign t[282] = t[327] ^ x[97];
  assign t[283] = t[328] ^ x[98];
  assign t[284] = t[329] ^ x[99];
  assign t[285] = t[330] ^ x[100];
  assign t[286] = t[331] ^ x[103];
  assign t[287] = t[332] ^ x[104];
  assign t[288] = t[333] ^ x[110];
  assign t[289] = t[334] ^ x[113];
  assign t[28] = x[7] ? t[46] : t[45];
  assign t[290] = t[335] ^ x[114];
  assign t[291] = t[336] ^ x[115];
  assign t[292] = t[337] ^ x[116];
  assign t[293] = t[338] ^ x[117];
  assign t[294] = t[339] ^ x[118];
  assign t[295] = t[340] ^ x[119];
  assign t[296] = t[341] ^ x[120];
  assign t[297] = t[342] ^ x[121];
  assign t[298] = t[343] ^ x[122];
  assign t[299] = t[344] ^ x[123];
  assign t[29] = x[7] ? t[48] : t[47];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[345] ^ x[124];
  assign t[301] = (~t[346] & t[347]);
  assign t[302] = (~t[348] & t[349]);
  assign t[303] = (~t[350] & t[351]);
  assign t[304] = (~t[352] & t[353]);
  assign t[305] = (~t[354] & t[355]);
  assign t[306] = (~t[356] & t[357]);
  assign t[307] = (~t[358] & t[359]);
  assign t[308] = (~t[356] & t[360]);
  assign t[309] = (~t[356] & t[361]);
  assign t[30] = ~(t[49]);
  assign t[310] = (~t[362] & t[363]);
  assign t[311] = (~t[364] & t[365]);
  assign t[312] = (~t[366] & t[367]);
  assign t[313] = (~t[358] & t[368]);
  assign t[314] = (~t[358] & t[369]);
  assign t[315] = (~t[370] & t[371]);
  assign t[316] = (~t[372] & t[373]);
  assign t[317] = (~t[374] & t[375]);
  assign t[318] = (~t[356] & t[376]);
  assign t[319] = (~t[362] & t[377]);
  assign t[31] = ~(t[50] | t[51]);
  assign t[320] = (~t[362] & t[378]);
  assign t[321] = (~t[364] & t[379]);
  assign t[322] = (~t[364] & t[380]);
  assign t[323] = (~t[366] & t[381]);
  assign t[324] = (~t[366] & t[382]);
  assign t[325] = (~t[383] & t[384]);
  assign t[326] = (~t[358] & t[385]);
  assign t[327] = (~t[370] & t[386]);
  assign t[328] = (~t[370] & t[387]);
  assign t[329] = (~t[372] & t[388]);
  assign t[32] = ~(t[52]);
  assign t[330] = (~t[372] & t[389]);
  assign t[331] = (~t[374] & t[390]);
  assign t[332] = (~t[374] & t[391]);
  assign t[333] = (~t[392] & t[393]);
  assign t[334] = (~t[362] & t[394]);
  assign t[335] = (~t[364] & t[395]);
  assign t[336] = (~t[366] & t[396]);
  assign t[337] = (~t[383] & t[397]);
  assign t[338] = (~t[383] & t[398]);
  assign t[339] = (~t[370] & t[399]);
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = (~t[372] & t[400]);
  assign t[341] = (~t[374] & t[401]);
  assign t[342] = (~t[392] & t[402]);
  assign t[343] = (~t[392] & t[403]);
  assign t[344] = (~t[383] & t[404]);
  assign t[345] = (~t[392] & t[405]);
  assign t[346] = t[406] ^ x[4];
  assign t[347] = t[407] ^ x[5];
  assign t[348] = t[408] ^ x[12];
  assign t[349] = t[409] ^ x[13];
  assign t[34] = ~(t[216] | t[55]);
  assign t[350] = t[410] ^ x[15];
  assign t[351] = t[411] ^ x[16];
  assign t[352] = t[412] ^ x[18];
  assign t[353] = t[413] ^ x[19];
  assign t[354] = t[414] ^ x[21];
  assign t[355] = t[415] ^ x[22];
  assign t[356] = t[416] ^ x[27];
  assign t[357] = t[417] ^ x[28];
  assign t[358] = t[418] ^ x[33];
  assign t[359] = t[419] ^ x[34];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[420] ^ x[35];
  assign t[361] = t[421] ^ x[36];
  assign t[362] = t[422] ^ x[41];
  assign t[363] = t[423] ^ x[42];
  assign t[364] = t[424] ^ x[49];
  assign t[365] = t[425] ^ x[50];
  assign t[366] = t[426] ^ x[55];
  assign t[367] = t[427] ^ x[56];
  assign t[368] = t[428] ^ x[57];
  assign t[369] = t[429] ^ x[58];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[430] ^ x[63];
  assign t[371] = t[431] ^ x[64];
  assign t[372] = t[432] ^ x[71];
  assign t[373] = t[433] ^ x[72];
  assign t[374] = t[434] ^ x[77];
  assign t[375] = t[435] ^ x[78];
  assign t[376] = t[436] ^ x[79];
  assign t[377] = t[437] ^ x[80];
  assign t[378] = t[438] ^ x[81];
  assign t[379] = t[439] ^ x[82];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[440] ^ x[83];
  assign t[381] = t[441] ^ x[86];
  assign t[382] = t[442] ^ x[87];
  assign t[383] = t[443] ^ x[92];
  assign t[384] = t[444] ^ x[93];
  assign t[385] = t[445] ^ x[96];
  assign t[386] = t[446] ^ x[97];
  assign t[387] = t[447] ^ x[98];
  assign t[388] = t[448] ^ x[99];
  assign t[389] = t[449] ^ x[100];
  assign t[38] = ~(t[47] ^ t[62]);
  assign t[390] = t[450] ^ x[103];
  assign t[391] = t[451] ^ x[104];
  assign t[392] = t[452] ^ x[109];
  assign t[393] = t[453] ^ x[110];
  assign t[394] = t[454] ^ x[113];
  assign t[395] = t[455] ^ x[114];
  assign t[396] = t[456] ^ x[115];
  assign t[397] = t[457] ^ x[116];
  assign t[398] = t[458] ^ x[117];
  assign t[399] = t[459] ^ x[118];
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[460] ^ x[119];
  assign t[401] = t[461] ^ x[120];
  assign t[402] = t[462] ^ x[121];
  assign t[403] = t[463] ^ x[122];
  assign t[404] = t[464] ^ x[123];
  assign t[405] = t[465] ^ x[124];
  assign t[406] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[407] = (x[0]);
  assign t[408] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[409] = (x[11]);
  assign t[40] = ~(t[65] ^ t[66]);
  assign t[410] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[411] = (x[14]);
  assign t[412] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[413] = (x[17]);
  assign t[414] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[415] = (x[20]);
  assign t[416] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[417] = (x[24]);
  assign t[418] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[419] = (x[30]);
  assign t[41] = ~(t[67] | t[68]);
  assign t[420] = (x[25]);
  assign t[421] = (x[26]);
  assign t[422] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[423] = (x[38]);
  assign t[424] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[425] = (x[46]);
  assign t[426] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[427] = (x[52]);
  assign t[428] = (x[31]);
  assign t[429] = (x[32]);
  assign t[42] = ~(t[217] | t[69]);
  assign t[430] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[431] = (x[60]);
  assign t[432] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[433] = (x[68]);
  assign t[434] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[435] = (x[74]);
  assign t[436] = (x[23]);
  assign t[437] = (x[39]);
  assign t[438] = (x[40]);
  assign t[439] = (x[47]);
  assign t[43] = ~(t[70] | t[71]);
  assign t[440] = (x[48]);
  assign t[441] = (x[53]);
  assign t[442] = (x[54]);
  assign t[443] = (x[88] & ~x[89] & ~x[90] & ~x[91]) | (~x[88] & x[89] & ~x[90] & ~x[91]) | (~x[88] & ~x[89] & x[90] & ~x[91]) | (~x[88] & ~x[89] & ~x[90] & x[91]) | (x[88] & x[89] & x[90] & ~x[91]) | (x[88] & x[89] & ~x[90] & x[91]) | (x[88] & ~x[89] & x[90] & x[91]) | (~x[88] & x[89] & x[90] & x[91]);
  assign t[444] = (x[89]);
  assign t[445] = (x[29]);
  assign t[446] = (x[61]);
  assign t[447] = (x[62]);
  assign t[448] = (x[69]);
  assign t[449] = (x[70]);
  assign t[44] = ~(t[72] ^ t[73]);
  assign t[450] = (x[75]);
  assign t[451] = (x[76]);
  assign t[452] = (x[105] & ~x[106] & ~x[107] & ~x[108]) | (~x[105] & x[106] & ~x[107] & ~x[108]) | (~x[105] & ~x[106] & x[107] & ~x[108]) | (~x[105] & ~x[106] & ~x[107] & x[108]) | (x[105] & x[106] & x[107] & ~x[108]) | (x[105] & x[106] & ~x[107] & x[108]) | (x[105] & ~x[106] & x[107] & x[108]) | (~x[105] & x[106] & x[107] & x[108]);
  assign t[453] = (x[106]);
  assign t[454] = (x[37]);
  assign t[455] = (x[45]);
  assign t[456] = (x[51]);
  assign t[457] = (x[90]);
  assign t[458] = (x[91]);
  assign t[459] = (x[59]);
  assign t[45] = ~(t[74] | t[75]);
  assign t[460] = (x[67]);
  assign t[461] = (x[73]);
  assign t[462] = (x[107]);
  assign t[463] = (x[108]);
  assign t[464] = (x[88]);
  assign t[465] = (x[105]);
  assign t[46] = ~(t[45] ^ t[76]);
  assign t[47] = ~(t[77] | t[78]);
  assign t[48] = ~(t[79] ^ t[80]);
  assign t[49] = ~(t[214]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[81] | t[82]);
  assign t[51] = ~(t[83] & t[84]);
  assign t[52] = ~(t[81] | t[85]);
  assign t[53] = ~(t[218]);
  assign t[54] = ~(t[219]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[220] | t[90]);
  assign t[58] = t[91] ? x[44] : x[43];
  assign t[59] = ~(t[92] & t[93]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[94] | t[95]);
  assign t[61] = ~(t[221] | t[96]);
  assign t[62] = ~(t[97] ^ t[98]);
  assign t[63] = ~(t[99] | t[100]);
  assign t[64] = ~(t[222] | t[101]);
  assign t[65] = ~(t[102] | t[103]);
  assign t[66] = ~(t[104] ^ t[105]);
  assign t[67] = ~(t[223]);
  assign t[68] = ~(t[224]);
  assign t[69] = ~(t[106] | t[107]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] | t[109]);
  assign t[71] = ~(t[225] | t[110]);
  assign t[72] = t[111] ? x[66] : x[65];
  assign t[73] = ~(t[112] & t[113]);
  assign t[74] = ~(t[114] | t[115]);
  assign t[75] = ~(t[226] | t[116]);
  assign t[76] = ~(t[117] ^ t[118]);
  assign t[77] = ~(t[119] | t[120]);
  assign t[78] = ~(t[227] | t[121]);
  assign t[79] = ~(t[122] | t[123]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[124] ^ t[125]);
  assign t[81] = ~(t[126]);
  assign t[82] = t[212] ? t[128] : t[127];
  assign t[83] = ~(t[129] | t[130]);
  assign t[84] = ~(t[131] | t[132]);
  assign t[85] = t[212] ? t[134] : t[133];
  assign t[86] = ~(t[228]);
  assign t[87] = ~(t[218] | t[219]);
  assign t[88] = ~(t[229]);
  assign t[89] = ~(t[230]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[135] | t[136]);
  assign t[91] = ~(t[49]);
  assign t[92] = ~(t[129] | t[137]);
  assign t[93] = ~(t[138] | t[139]);
  assign t[94] = ~(t[231]);
  assign t[95] = ~(t[232]);
  assign t[96] = ~(t[140] | t[141]);
  assign t[97] = t[91] ? x[85] : x[84];
  assign t[98] = ~(t[142] & t[143]);
  assign t[99] = ~(t[233]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [163:0] x;
 output y;

 wire [634:0] t;
  assign t[0] = t[1] ? t[2] : t[387];
  assign t[100] = ~(t[409]);
  assign t[101] = ~(t[398] | t[399]);
  assign t[102] = ~(t[410]);
  assign t[103] = ~(t[411]);
  assign t[104] = ~(t[140] | t[141]);
  assign t[105] = ~(t[48]);
  assign t[106] = ~(t[129] | t[142]);
  assign t[107] = ~(t[127]);
  assign t[108] = ~(t[412]);
  assign t[109] = ~(t[413]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[143] | t[144]);
  assign t[111] = t[30] ? x[94] : x[93];
  assign t[112] = ~(t[145] & t[146]);
  assign t[113] = ~(t[414]);
  assign t[114] = ~(t[415]);
  assign t[115] = ~(t[147] | t[148]);
  assign t[116] = ~(t[149] | t[150]);
  assign t[117] = ~(t[416] | t[151]);
  assign t[118] = t[30] ? x[104] : x[103];
  assign t[119] = ~(t[83] & t[152]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[390]);
  assign t[121] = ~(t[391] & t[153]);
  assign t[122] = ~(x[7] & t[154]);
  assign t[123] = ~(t[155] & t[391]);
  assign t[124] = ~(t[156] & t[157]);
  assign t[125] = ~(t[120] | t[158]);
  assign t[126] = ~(t[120] | t[159]);
  assign t[127] = ~(t[79] | t[160]);
  assign t[128] = ~(t[161] & t[162]);
  assign t[129] = ~(t[79] | t[163]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[417]);
  assign t[131] = ~(t[404] | t[405]);
  assign t[132] = ~(t[418]);
  assign t[133] = ~(t[419]);
  assign t[134] = ~(t[164] | t[165]);
  assign t[135] = ~(t[138] | t[166]);
  assign t[136] = ~(t[420]);
  assign t[137] = ~(t[407] | t[408]);
  assign t[138] = ~(t[167] & t[168]);
  assign t[139] = ~(t[169] & t[31]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[421]);
  assign t[141] = ~(t[410] | t[411]);
  assign t[142] = ~(t[170] & t[83]);
  assign t[143] = ~(t[422]);
  assign t[144] = ~(t[412] | t[413]);
  assign t[145] = ~(t[171] | t[126]);
  assign t[146] = ~(t[172] | t[173]);
  assign t[147] = ~(t[423]);
  assign t[148] = ~(t[414] | t[415]);
  assign t[149] = ~(t[424]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[425]);
  assign t[151] = ~(t[174] | t[175]);
  assign t[152] = ~(t[176] | t[177]);
  assign t[153] = ~(x[7] | t[178]);
  assign t[154] = ~(t[389] | t[391]);
  assign t[155] = ~(x[7] | t[389]);
  assign t[156] = x[7] & t[389];
  assign t[157] = ~(t[391]);
  assign t[158] = t[388] ? t[124] : t[179];
  assign t[159] = t[388] ? t[180] : t[122];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[388] ? t[179] : t[181];
  assign t[161] = ~(t[182] | t[49]);
  assign t[162] = ~(t[51] & t[183]);
  assign t[163] = t[388] ? t[184] : t[180];
  assign t[164] = ~(t[426]);
  assign t[165] = ~(t[418] | t[419]);
  assign t[166] = ~(t[185] & t[186]);
  assign t[167] = ~(t[82] & t[187]);
  assign t[168] = ~(t[188] & t[189]);
  assign t[169] = ~(t[127] | t[190]);
  assign t[16] = ~(t[388] & t[389]);
  assign t[170] = ~(t[182] | t[176]);
  assign t[171] = ~(t[120] | t[191]);
  assign t[172] = ~(t[87]);
  assign t[173] = ~(t[79] | t[192]);
  assign t[174] = ~(t[427]);
  assign t[175] = ~(t[424] | t[425]);
  assign t[176] = ~(t[193] & t[194]);
  assign t[177] = ~(t[162] & t[186]);
  assign t[178] = ~(t[389]);
  assign t[179] = ~(t[155] & t[157]);
  assign t[17] = ~(t[390] & t[391]);
  assign t[180] = ~(t[153] & t[157]);
  assign t[181] = ~(t[156] & t[391]);
  assign t[182] = ~(t[79] | t[195]);
  assign t[183] = t[155] | t[156];
  assign t[184] = ~(x[7] & t[188]);
  assign t[185] = ~(t[126]);
  assign t[186] = t[120] | t[196];
  assign t[187] = ~(t[121] & t[184]);
  assign t[188] = ~(t[389] | t[157]);
  assign t[189] = t[79] & t[388];
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[79] | t[197]);
  assign t[191] = t[388] ? t[179] : t[124];
  assign t[192] = t[388] ? t[121] : t[122];
  assign t[193] = ~(t[171] | t[198]);
  assign t[194] = ~(t[120] & t[199]);
  assign t[195] = t[388] ? t[181] : t[179];
  assign t[196] = t[388] ? t[122] : t[180];
  assign t[197] = t[388] ? t[123] : t[124];
  assign t[198] = ~(t[79] | t[200]);
  assign t[199] = ~(t[122] & t[121]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[388] ? t[180] : t[184];
  assign t[201] = t[1] ? t[202] : t[428];
  assign t[202] = x[6] ? t[204] : t[203];
  assign t[203] = x[7] ? t[206] : t[205];
  assign t[204] = t[207] ^ x[117];
  assign t[205] = t[208] ^ t[209];
  assign t[206] = ~(t[210] ^ t[211]);
  assign t[207] = x[118] ^ x[119];
  assign t[208] = t[30] ? x[119] : x[118];
  assign t[209] = ~(t[212] ^ t[213]);
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = x[7] ? t[215] : t[214];
  assign t[211] = ~(t[216] ^ t[217]);
  assign t[212] = x[7] ? t[219] : t[218];
  assign t[213] = ~(t[220] ^ t[221]);
  assign t[214] = ~(t[222] & t[223]);
  assign t[215] = t[224] ^ t[218];
  assign t[216] = x[7] ? t[226] : t[225];
  assign t[217] = x[7] ? t[228] : t[227];
  assign t[218] = ~(t[229] & t[230]);
  assign t[219] = t[231] ^ t[232];
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = x[7] ? t[234] : t[233];
  assign t[221] = x[7] ? t[236] : t[235];
  assign t[222] = ~(t[394] & t[54]);
  assign t[223] = ~(t[403] & t[237]);
  assign t[224] = t[390] ? x[121] : x[120];
  assign t[225] = ~(t[238] & t[239]);
  assign t[226] = t[240] ^ t[225];
  assign t[227] = ~(t[241] & t[242]);
  assign t[228] = t[243] ^ t[244];
  assign t[229] = ~(t[398] & t[66]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = ~(t[409] & t[245]);
  assign t[231] = t[105] ? x[123] : x[122];
  assign t[232] = ~(t[246] & t[247]);
  assign t[233] = ~(t[248] & t[249]);
  assign t[234] = t[250] ^ t[251];
  assign t[235] = ~(t[252] & t[253]);
  assign t[236] = t[254] ^ t[235];
  assign t[237] = ~(t[395] & t[53]);
  assign t[238] = ~(t[407] & t[96]);
  assign t[239] = ~(t[420] & t[255]);
  assign t[23] = ~(t[26] ^ t[35]);
  assign t[240] = t[390] ? x[125] : x[124];
  assign t[241] = ~(t[404] & t[89]);
  assign t[242] = ~(t[417] & t[256]);
  assign t[243] = t[390] ? x[127] : x[126];
  assign t[244] = ~(t[257] & t[258]);
  assign t[245] = ~(t[399] & t[65]);
  assign t[246] = ~(t[410] & t[103]);
  assign t[247] = ~(t[421] & t[259]);
  assign t[248] = ~(t[414] & t[114]);
  assign t[249] = ~(t[423] & t[260]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[30] ? x[129] : x[128];
  assign t[251] = ~(t[261] & t[262]);
  assign t[252] = ~(t[412] & t[109]);
  assign t[253] = ~(t[422] & t[263]);
  assign t[254] = t[30] ? x[131] : x[130];
  assign t[255] = ~(t[408] & t[95]);
  assign t[256] = ~(t[405] & t[88]);
  assign t[257] = ~(t[418] & t[133]);
  assign t[258] = ~(t[426] & t[264]);
  assign t[259] = ~(t[411] & t[102]);
  assign t[25] = x[7] ? t[39] : t[38];
  assign t[260] = ~(t[415] & t[113]);
  assign t[261] = ~(t[424] & t[150]);
  assign t[262] = ~(t[427] & t[265]);
  assign t[263] = ~(t[413] & t[108]);
  assign t[264] = ~(t[419] & t[132]);
  assign t[265] = ~(t[425] & t[149]);
  assign t[266] = t[1] ? t[267] : t[429];
  assign t[267] = x[6] ? t[269] : t[268];
  assign t[268] = x[7] ? t[271] : t[270];
  assign t[269] = t[272] ^ x[133];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[273] ^ t[274];
  assign t[271] = ~(t[275] ^ t[276]);
  assign t[272] = x[134] ^ x[135];
  assign t[273] = t[30] ? x[135] : x[134];
  assign t[274] = ~(t[277] ^ t[278]);
  assign t[275] = x[7] ? t[280] : t[279];
  assign t[276] = ~(t[281] ^ t[282]);
  assign t[277] = x[7] ? t[284] : t[283];
  assign t[278] = ~(t[285] ^ t[286]);
  assign t[279] = ~(t[287] & t[288]);
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[289] ^ t[283];
  assign t[281] = x[7] ? t[291] : t[290];
  assign t[282] = x[7] ? t[293] : t[292];
  assign t[283] = ~(t[294] & t[295]);
  assign t[284] = t[296] ^ t[297];
  assign t[285] = x[7] ? t[299] : t[298];
  assign t[286] = x[7] ? t[301] : t[300];
  assign t[287] = ~(t[54] & t[84]);
  assign t[288] = ~(t[302] & t[392]);
  assign t[289] = t[390] ? x[137] : x[136];
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = ~(t[303] & t[304]);
  assign t[291] = t[305] ^ t[306];
  assign t[292] = ~(t[307] & t[308]);
  assign t[293] = t[309] ^ t[292];
  assign t[294] = ~(t[66] & t[100]);
  assign t[295] = ~(t[310] & t[393]);
  assign t[296] = t[105] ? x[139] : x[138];
  assign t[297] = ~(t[311] & t[312]);
  assign t[298] = ~(t[313] & t[314]);
  assign t[299] = t[315] ^ t[298];
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = ~(t[316] & t[317]);
  assign t[301] = t[318] ^ t[319];
  assign t[302] = ~(t[320] & t[53]);
  assign t[303] = ~(t[89] & t[130]);
  assign t[304] = ~(t[321] & t[396]);
  assign t[305] = t[390] ? x[141] : x[140];
  assign t[306] = ~(t[322] & t[323]);
  assign t[307] = ~(t[96] & t[136]);
  assign t[308] = ~(t[324] & t[397]);
  assign t[309] = t[390] ? x[143] : x[142];
  assign t[30] = ~(t[48]);
  assign t[310] = ~(t[325] & t[65]);
  assign t[311] = ~(t[103] & t[140]);
  assign t[312] = ~(t[326] & t[400]);
  assign t[313] = ~(t[109] & t[143]);
  assign t[314] = ~(t[327] & t[401]);
  assign t[315] = t[30] ? x[145] : x[144];
  assign t[316] = ~(t[114] & t[147]);
  assign t[317] = ~(t[328] & t[402]);
  assign t[318] = t[30] ? x[147] : x[146];
  assign t[319] = ~(t[329] & t[330]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = ~(t[403] & t[395]);
  assign t[321] = ~(t[331] & t[88]);
  assign t[322] = ~(t[133] & t[164]);
  assign t[323] = ~(t[332] & t[406]);
  assign t[324] = ~(t[333] & t[95]);
  assign t[325] = ~(t[409] & t[399]);
  assign t[326] = ~(t[334] & t[102]);
  assign t[327] = ~(t[335] & t[108]);
  assign t[328] = ~(t[336] & t[113]);
  assign t[329] = ~(t[150] & t[174]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = ~(t[337] & t[416]);
  assign t[331] = ~(t[417] & t[405]);
  assign t[332] = ~(t[338] & t[132]);
  assign t[333] = ~(t[420] & t[408]);
  assign t[334] = ~(t[421] & t[411]);
  assign t[335] = ~(t[422] & t[413]);
  assign t[336] = ~(t[423] & t[415]);
  assign t[337] = ~(t[339] & t[149]);
  assign t[338] = ~(t[426] & t[419]);
  assign t[339] = ~(t[427] & t[425]);
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[1] ? t[341] : t[430];
  assign t[341] = x[6] ? t[343] : t[342];
  assign t[342] = x[7] ? t[345] : t[344];
  assign t[343] = t[346] ^ x[149];
  assign t[344] = t[347] ^ t[348];
  assign t[345] = ~(t[349] ^ t[350]);
  assign t[346] = x[150] ^ x[151];
  assign t[347] = t[30] ? x[151] : x[150];
  assign t[348] = ~(t[351] ^ t[352]);
  assign t[349] = x[7] ? t[354] : t[353];
  assign t[34] = ~(t[392] | t[55]);
  assign t[350] = ~(t[355] ^ t[356]);
  assign t[351] = x[7] ? t[358] : t[357];
  assign t[352] = ~(t[359] ^ t[360]);
  assign t[353] = ~(t[287] & t[361]);
  assign t[354] = t[362] ^ t[357];
  assign t[355] = x[7] ? t[364] : t[363];
  assign t[356] = x[7] ? t[366] : t[365];
  assign t[357] = ~(t[294] & t[367]);
  assign t[358] = t[368] ^ t[369];
  assign t[359] = x[7] ? t[371] : t[370];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = x[7] ? t[373] : t[372];
  assign t[361] = t[33] | t[392];
  assign t[362] = t[390] ? x[153] : x[152];
  assign t[363] = ~(t[303] & t[374]);
  assign t[364] = t[375] ^ t[376];
  assign t[365] = ~(t[307] & t[377]);
  assign t[366] = t[378] ^ t[365];
  assign t[367] = t[40] | t[393];
  assign t[368] = t[105] ? x[155] : x[154];
  assign t[369] = ~(t[311] & t[379]);
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = ~(t[313] & t[380]);
  assign t[371] = t[381] ^ t[370];
  assign t[372] = ~(t[316] & t[382]);
  assign t[373] = t[383] ^ t[384];
  assign t[374] = t[58] | t[396];
  assign t[375] = t[390] ? x[157] : x[156];
  assign t[376] = ~(t[322] & t[385]);
  assign t[377] = t[62] | t[397];
  assign t[378] = t[390] ? x[159] : x[158];
  assign t[379] = t[68] | t[400];
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[380] = t[72] | t[401];
  assign t[381] = t[30] ? x[161] : x[160];
  assign t[382] = t[75] | t[402];
  assign t[383] = t[30] ? x[163] : x[162];
  assign t[384] = ~(t[329] & t[386]);
  assign t[385] = t[91] | t[406];
  assign t[386] = t[116] | t[416];
  assign t[387] = (t[431]);
  assign t[388] = (t[432]);
  assign t[389] = (t[433]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[390] = (t[434]);
  assign t[391] = (t[435]);
  assign t[392] = (t[436]);
  assign t[393] = (t[437]);
  assign t[394] = (t[438]);
  assign t[395] = (t[439]);
  assign t[396] = (t[440]);
  assign t[397] = (t[441]);
  assign t[398] = (t[442]);
  assign t[399] = (t[443]);
  assign t[39] = ~(t[38] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (t[444]);
  assign t[401] = (t[445]);
  assign t[402] = (t[446]);
  assign t[403] = (t[447]);
  assign t[404] = (t[448]);
  assign t[405] = (t[449]);
  assign t[406] = (t[450]);
  assign t[407] = (t[451]);
  assign t[408] = (t[452]);
  assign t[409] = (t[453]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (t[454]);
  assign t[411] = (t[455]);
  assign t[412] = (t[456]);
  assign t[413] = (t[457]);
  assign t[414] = (t[458]);
  assign t[415] = (t[459]);
  assign t[416] = (t[460]);
  assign t[417] = (t[461]);
  assign t[418] = (t[462]);
  assign t[419] = (t[463]);
  assign t[41] = ~(t[393] | t[67]);
  assign t[420] = (t[464]);
  assign t[421] = (t[465]);
  assign t[422] = (t[466]);
  assign t[423] = (t[467]);
  assign t[424] = (t[468]);
  assign t[425] = (t[469]);
  assign t[426] = (t[470]);
  assign t[427] = (t[471]);
  assign t[428] = (t[472]);
  assign t[429] = (t[473]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (t[474]);
  assign t[431] = t[475] ^ x[5];
  assign t[432] = t[476] ^ x[13];
  assign t[433] = t[477] ^ x[16];
  assign t[434] = t[478] ^ x[19];
  assign t[435] = t[479] ^ x[22];
  assign t[436] = t[480] ^ x[28];
  assign t[437] = t[481] ^ x[34];
  assign t[438] = t[482] ^ x[35];
  assign t[439] = t[483] ^ x[36];
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[440] = t[484] ^ x[44];
  assign t[441] = t[485] ^ x[50];
  assign t[442] = t[486] ^ x[51];
  assign t[443] = t[487] ^ x[52];
  assign t[444] = t[488] ^ x[58];
  assign t[445] = t[489] ^ x[66];
  assign t[446] = t[490] ^ x[72];
  assign t[447] = t[491] ^ x[73];
  assign t[448] = t[492] ^ x[74];
  assign t[449] = t[493] ^ x[75];
  assign t[44] = ~(t[72] | t[73]);
  assign t[450] = t[494] ^ x[81];
  assign t[451] = t[495] ^ x[84];
  assign t[452] = t[496] ^ x[85];
  assign t[453] = t[497] ^ x[88];
  assign t[454] = t[498] ^ x[89];
  assign t[455] = t[499] ^ x[90];
  assign t[456] = t[500] ^ x[91];
  assign t[457] = t[501] ^ x[92];
  assign t[458] = t[502] ^ x[95];
  assign t[459] = t[503] ^ x[96];
  assign t[45] = ~(t[44] ^ t[74]);
  assign t[460] = t[504] ^ x[102];
  assign t[461] = t[505] ^ x[105];
  assign t[462] = t[506] ^ x[106];
  assign t[463] = t[507] ^ x[107];
  assign t[464] = t[508] ^ x[108];
  assign t[465] = t[509] ^ x[109];
  assign t[466] = t[510] ^ x[110];
  assign t[467] = t[511] ^ x[111];
  assign t[468] = t[512] ^ x[112];
  assign t[469] = t[513] ^ x[113];
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = t[514] ^ x[114];
  assign t[471] = t[515] ^ x[115];
  assign t[472] = t[516] ^ x[116];
  assign t[473] = t[517] ^ x[132];
  assign t[474] = t[518] ^ x[148];
  assign t[475] = (~t[519] & t[520]);
  assign t[476] = (~t[521] & t[522]);
  assign t[477] = (~t[523] & t[524]);
  assign t[478] = (~t[525] & t[526]);
  assign t[479] = (~t[527] & t[528]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (~t[529] & t[530]);
  assign t[481] = (~t[531] & t[532]);
  assign t[482] = (~t[529] & t[533]);
  assign t[483] = (~t[529] & t[534]);
  assign t[484] = (~t[535] & t[536]);
  assign t[485] = (~t[537] & t[538]);
  assign t[486] = (~t[531] & t[539]);
  assign t[487] = (~t[531] & t[540]);
  assign t[488] = (~t[541] & t[542]);
  assign t[489] = (~t[543] & t[544]);
  assign t[48] = ~(t[390]);
  assign t[490] = (~t[545] & t[546]);
  assign t[491] = (~t[529] & t[547]);
  assign t[492] = (~t[535] & t[548]);
  assign t[493] = (~t[535] & t[549]);
  assign t[494] = (~t[550] & t[551]);
  assign t[495] = (~t[537] & t[552]);
  assign t[496] = (~t[537] & t[553]);
  assign t[497] = (~t[531] & t[554]);
  assign t[498] = (~t[541] & t[555]);
  assign t[499] = (~t[541] & t[556]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[543] & t[557]);
  assign t[501] = (~t[543] & t[558]);
  assign t[502] = (~t[545] & t[559]);
  assign t[503] = (~t[545] & t[560]);
  assign t[504] = (~t[561] & t[562]);
  assign t[505] = (~t[535] & t[563]);
  assign t[506] = (~t[550] & t[564]);
  assign t[507] = (~t[550] & t[565]);
  assign t[508] = (~t[537] & t[566]);
  assign t[509] = (~t[541] & t[567]);
  assign t[50] = ~(t[79] | t[81]);
  assign t[510] = (~t[543] & t[568]);
  assign t[511] = (~t[545] & t[569]);
  assign t[512] = (~t[561] & t[570]);
  assign t[513] = (~t[561] & t[571]);
  assign t[514] = (~t[550] & t[572]);
  assign t[515] = (~t[561] & t[573]);
  assign t[516] = (~t[519] & t[574]);
  assign t[517] = (~t[519] & t[575]);
  assign t[518] = (~t[519] & t[576]);
  assign t[519] = t[577] ^ x[4];
  assign t[51] = t[391] & t[82];
  assign t[520] = t[578] ^ x[5];
  assign t[521] = t[579] ^ x[12];
  assign t[522] = t[580] ^ x[13];
  assign t[523] = t[581] ^ x[15];
  assign t[524] = t[582] ^ x[16];
  assign t[525] = t[583] ^ x[18];
  assign t[526] = t[584] ^ x[19];
  assign t[527] = t[585] ^ x[21];
  assign t[528] = t[586] ^ x[22];
  assign t[529] = t[587] ^ x[27];
  assign t[52] = ~(t[83]);
  assign t[530] = t[588] ^ x[28];
  assign t[531] = t[589] ^ x[33];
  assign t[532] = t[590] ^ x[34];
  assign t[533] = t[591] ^ x[35];
  assign t[534] = t[592] ^ x[36];
  assign t[535] = t[593] ^ x[43];
  assign t[536] = t[594] ^ x[44];
  assign t[537] = t[595] ^ x[49];
  assign t[538] = t[596] ^ x[50];
  assign t[539] = t[597] ^ x[51];
  assign t[53] = ~(t[394]);
  assign t[540] = t[598] ^ x[52];
  assign t[541] = t[599] ^ x[57];
  assign t[542] = t[600] ^ x[58];
  assign t[543] = t[601] ^ x[65];
  assign t[544] = t[602] ^ x[66];
  assign t[545] = t[603] ^ x[71];
  assign t[546] = t[604] ^ x[72];
  assign t[547] = t[605] ^ x[73];
  assign t[548] = t[606] ^ x[74];
  assign t[549] = t[607] ^ x[75];
  assign t[54] = ~(t[395]);
  assign t[550] = t[608] ^ x[80];
  assign t[551] = t[609] ^ x[81];
  assign t[552] = t[610] ^ x[84];
  assign t[553] = t[611] ^ x[85];
  assign t[554] = t[612] ^ x[88];
  assign t[555] = t[613] ^ x[89];
  assign t[556] = t[614] ^ x[90];
  assign t[557] = t[615] ^ x[91];
  assign t[558] = t[616] ^ x[92];
  assign t[559] = t[617] ^ x[95];
  assign t[55] = ~(t[84] | t[85]);
  assign t[560] = t[618] ^ x[96];
  assign t[561] = t[619] ^ x[101];
  assign t[562] = t[620] ^ x[102];
  assign t[563] = t[621] ^ x[105];
  assign t[564] = t[622] ^ x[106];
  assign t[565] = t[623] ^ x[107];
  assign t[566] = t[624] ^ x[108];
  assign t[567] = t[625] ^ x[109];
  assign t[568] = t[626] ^ x[110];
  assign t[569] = t[627] ^ x[111];
  assign t[56] = t[390] ? x[38] : x[37];
  assign t[570] = t[628] ^ x[112];
  assign t[571] = t[629] ^ x[113];
  assign t[572] = t[630] ^ x[114];
  assign t[573] = t[631] ^ x[115];
  assign t[574] = t[632] ^ x[116];
  assign t[575] = t[633] ^ x[132];
  assign t[576] = t[634] ^ x[148];
  assign t[577] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[578] = (x[0]);
  assign t[579] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = ~(t[86] & t[87]);
  assign t[580] = (x[11]);
  assign t[581] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[582] = (x[14]);
  assign t[583] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[584] = (x[17]);
  assign t[585] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[586] = (x[20]);
  assign t[587] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[588] = (x[24]);
  assign t[589] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[58] = ~(t[88] | t[89]);
  assign t[590] = (x[30]);
  assign t[591] = (x[25]);
  assign t[592] = (x[26]);
  assign t[593] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[594] = (x[40]);
  assign t[595] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[596] = (x[46]);
  assign t[597] = (x[31]);
  assign t[598] = (x[32]);
  assign t[599] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[59] = ~(t[396] | t[90]);
  assign t[5] = t[9] ^ x[8];
  assign t[600] = (x[54]);
  assign t[601] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[602] = (x[62]);
  assign t[603] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[604] = (x[68]);
  assign t[605] = (x[23]);
  assign t[606] = (x[41]);
  assign t[607] = (x[42]);
  assign t[608] = (x[76] & ~x[77] & ~x[78] & ~x[79]) | (~x[76] & x[77] & ~x[78] & ~x[79]) | (~x[76] & ~x[77] & x[78] & ~x[79]) | (~x[76] & ~x[77] & ~x[78] & x[79]) | (x[76] & x[77] & x[78] & ~x[79]) | (x[76] & x[77] & ~x[78] & x[79]) | (x[76] & ~x[77] & x[78] & x[79]) | (~x[76] & x[77] & x[78] & x[79]);
  assign t[609] = (x[77]);
  assign t[60] = ~(t[91] | t[92]);
  assign t[610] = (x[47]);
  assign t[611] = (x[48]);
  assign t[612] = (x[29]);
  assign t[613] = (x[55]);
  assign t[614] = (x[56]);
  assign t[615] = (x[63]);
  assign t[616] = (x[64]);
  assign t[617] = (x[69]);
  assign t[618] = (x[70]);
  assign t[619] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[61] = ~(t[93] ^ t[94]);
  assign t[620] = (x[98]);
  assign t[621] = (x[39]);
  assign t[622] = (x[78]);
  assign t[623] = (x[79]);
  assign t[624] = (x[45]);
  assign t[625] = (x[53]);
  assign t[626] = (x[61]);
  assign t[627] = (x[67]);
  assign t[628] = (x[99]);
  assign t[629] = (x[100]);
  assign t[62] = ~(t[95] | t[96]);
  assign t[630] = (x[76]);
  assign t[631] = (x[97]);
  assign t[632] = (x[1]);
  assign t[633] = (x[2]);
  assign t[634] = (x[3]);
  assign t[63] = ~(t[397] | t[97]);
  assign t[64] = ~(t[98] ^ t[99]);
  assign t[65] = ~(t[398]);
  assign t[66] = ~(t[399]);
  assign t[67] = ~(t[100] | t[101]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[400] | t[104]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[105] ? x[60] : x[59];
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[108] | t[109]);
  assign t[73] = ~(t[401] | t[110]);
  assign t[74] = ~(t[111] ^ t[112]);
  assign t[75] = ~(t[113] | t[114]);
  assign t[76] = ~(t[402] | t[115]);
  assign t[77] = ~(t[116] | t[117]);
  assign t[78] = ~(t[118] ^ t[119]);
  assign t[79] = ~(t[120]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[388] ? t[122] : t[121];
  assign t[81] = t[388] ? t[124] : t[123];
  assign t[82] = ~(t[120] | t[388]);
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = ~(t[403]);
  assign t[85] = ~(t[394] | t[395]);
  assign t[86] = ~(t[127] | t[128]);
  assign t[87] = ~(t[129] | t[50]);
  assign t[88] = ~(t[404]);
  assign t[89] = ~(t[405]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[130] | t[131]);
  assign t[91] = ~(t[132] | t[133]);
  assign t[92] = ~(t[406] | t[134]);
  assign t[93] = t[105] ? x[83] : x[82];
  assign t[94] = ~(t[135] & t[107]);
  assign t[95] = ~(t[407]);
  assign t[96] = ~(t[408]);
  assign t[97] = ~(t[136] | t[137]);
  assign t[98] = t[390] ? x[87] : x[86];
  assign t[99] = t[138] | t[139];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[201] & ~t[266] & ~t[340]) | (~t[0] & t[201] & ~t[266] & ~t[340]) | (~t[0] & ~t[201] & t[266] & ~t[340]) | (~t[0] & ~t[201] & ~t[266] & t[340]) | (t[0] & t[201] & t[266] & ~t[340]) | (t[0] & t[201] & ~t[266] & t[340]) | (t[0] & ~t[201] & t[266] & t[340]) | (~t[0] & t[201] & t[266] & t[340]);
endmodule

module R2ind176(x, y);
 input [115:0] x;
 output y;

 wire [334:0] t;
  assign t[0] = t[1] ? t[2] : t[102];
  assign t[100] = ~(t[141]);
  assign t[101] = ~(t[142]);
  assign t[102] = (t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = t[184] ^ x[5];
  assign t[144] = t[185] ^ x[13];
  assign t[145] = t[186] ^ x[16];
  assign t[146] = t[187] ^ x[19];
  assign t[147] = t[188] ^ x[22];
  assign t[148] = t[189] ^ x[28];
  assign t[149] = t[190] ^ x[36];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[39];
  assign t[151] = t[192] ^ x[40];
  assign t[152] = t[193] ^ x[46];
  assign t[153] = t[194] ^ x[54];
  assign t[154] = t[195] ^ x[57];
  assign t[155] = t[196] ^ x[58];
  assign t[156] = t[197] ^ x[64];
  assign t[157] = t[198] ^ x[70];
  assign t[158] = t[199] ^ x[78];
  assign t[159] = t[200] ^ x[81];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[82];
  assign t[161] = t[202] ^ x[83];
  assign t[162] = t[203] ^ x[89];
  assign t[163] = t[204] ^ x[90];
  assign t[164] = t[205] ^ x[91];
  assign t[165] = t[206] ^ x[92];
  assign t[166] = t[207] ^ x[93];
  assign t[167] = t[208] ^ x[94];
  assign t[168] = t[209] ^ x[95];
  assign t[169] = t[210] ^ x[96];
  assign t[16] = ~(t[103] & t[104]);
  assign t[170] = t[211] ^ x[97];
  assign t[171] = t[212] ^ x[98];
  assign t[172] = t[213] ^ x[104];
  assign t[173] = t[214] ^ x[105];
  assign t[174] = t[215] ^ x[106];
  assign t[175] = t[216] ^ x[107];
  assign t[176] = t[217] ^ x[108];
  assign t[177] = t[218] ^ x[109];
  assign t[178] = t[219] ^ x[110];
  assign t[179] = t[220] ^ x[111];
  assign t[17] = ~(t[105] & t[106]);
  assign t[180] = t[221] ^ x[112];
  assign t[181] = t[222] ^ x[113];
  assign t[182] = t[223] ^ x[114];
  assign t[183] = t[224] ^ x[115];
  assign t[184] = (~t[225] & t[226]);
  assign t[185] = (~t[227] & t[228]);
  assign t[186] = (~t[229] & t[230]);
  assign t[187] = (~t[231] & t[232]);
  assign t[188] = (~t[233] & t[234]);
  assign t[189] = (~t[235] & t[236]);
  assign t[18] = ~(t[25]);
  assign t[190] = (~t[237] & t[238]);
  assign t[191] = (~t[235] & t[239]);
  assign t[192] = (~t[235] & t[240]);
  assign t[193] = (~t[241] & t[242]);
  assign t[194] = (~t[243] & t[244]);
  assign t[195] = (~t[237] & t[245]);
  assign t[196] = (~t[237] & t[246]);
  assign t[197] = (~t[247] & t[248]);
  assign t[198] = (~t[249] & t[250]);
  assign t[199] = (~t[251] & t[252]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[235] & t[253]);
  assign t[201] = (~t[241] & t[254]);
  assign t[202] = (~t[241] & t[255]);
  assign t[203] = (~t[256] & t[257]);
  assign t[204] = (~t[243] & t[258]);
  assign t[205] = (~t[243] & t[259]);
  assign t[206] = (~t[237] & t[260]);
  assign t[207] = (~t[247] & t[261]);
  assign t[208] = (~t[247] & t[262]);
  assign t[209] = (~t[249] & t[263]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[249] & t[264]);
  assign t[211] = (~t[251] & t[265]);
  assign t[212] = (~t[251] & t[266]);
  assign t[213] = (~t[267] & t[268]);
  assign t[214] = (~t[241] & t[269]);
  assign t[215] = (~t[256] & t[270]);
  assign t[216] = (~t[256] & t[271]);
  assign t[217] = (~t[243] & t[272]);
  assign t[218] = (~t[247] & t[273]);
  assign t[219] = (~t[249] & t[274]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[251] & t[275]);
  assign t[221] = (~t[267] & t[276]);
  assign t[222] = (~t[267] & t[277]);
  assign t[223] = (~t[256] & t[278]);
  assign t[224] = (~t[267] & t[279]);
  assign t[225] = t[280] ^ x[4];
  assign t[226] = t[281] ^ x[5];
  assign t[227] = t[282] ^ x[12];
  assign t[228] = t[283] ^ x[13];
  assign t[229] = t[284] ^ x[15];
  assign t[22] = t[32] ^ t[26];
  assign t[230] = t[285] ^ x[16];
  assign t[231] = t[286] ^ x[18];
  assign t[232] = t[287] ^ x[19];
  assign t[233] = t[288] ^ x[21];
  assign t[234] = t[289] ^ x[22];
  assign t[235] = t[290] ^ x[27];
  assign t[236] = t[291] ^ x[28];
  assign t[237] = t[292] ^ x[35];
  assign t[238] = t[293] ^ x[36];
  assign t[239] = t[294] ^ x[39];
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = t[295] ^ x[40];
  assign t[241] = t[296] ^ x[45];
  assign t[242] = t[297] ^ x[46];
  assign t[243] = t[298] ^ x[53];
  assign t[244] = t[299] ^ x[54];
  assign t[245] = t[300] ^ x[57];
  assign t[246] = t[301] ^ x[58];
  assign t[247] = t[302] ^ x[63];
  assign t[248] = t[303] ^ x[64];
  assign t[249] = t[304] ^ x[69];
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = t[305] ^ x[70];
  assign t[251] = t[306] ^ x[77];
  assign t[252] = t[307] ^ x[78];
  assign t[253] = t[308] ^ x[81];
  assign t[254] = t[309] ^ x[82];
  assign t[255] = t[310] ^ x[83];
  assign t[256] = t[311] ^ x[88];
  assign t[257] = t[312] ^ x[89];
  assign t[258] = t[313] ^ x[90];
  assign t[259] = t[314] ^ x[91];
  assign t[25] = ~(t[105]);
  assign t[260] = t[315] ^ x[92];
  assign t[261] = t[316] ^ x[93];
  assign t[262] = t[317] ^ x[94];
  assign t[263] = t[318] ^ x[95];
  assign t[264] = t[319] ^ x[96];
  assign t[265] = t[320] ^ x[97];
  assign t[266] = t[321] ^ x[98];
  assign t[267] = t[322] ^ x[103];
  assign t[268] = t[323] ^ x[104];
  assign t[269] = t[324] ^ x[105];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[325] ^ x[106];
  assign t[271] = t[326] ^ x[107];
  assign t[272] = t[327] ^ x[108];
  assign t[273] = t[328] ^ x[109];
  assign t[274] = t[329] ^ x[110];
  assign t[275] = t[330] ^ x[111];
  assign t[276] = t[331] ^ x[112];
  assign t[277] = t[332] ^ x[113];
  assign t[278] = t[333] ^ x[114];
  assign t[279] = t[334] ^ x[115];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[281] = (x[3]);
  assign t[282] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[283] = (x[11]);
  assign t[284] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[285] = (x[14]);
  assign t[286] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[287] = (x[17]);
  assign t[288] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[289] = (x[20]);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[290] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[291] = (x[24]);
  assign t[292] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[293] = (x[32]);
  assign t[294] = (x[26]);
  assign t[295] = (x[23]);
  assign t[296] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[297] = (x[42]);
  assign t[298] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[299] = (x[50]);
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[34]);
  assign t[301] = (x[31]);
  assign t[302] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[303] = (x[60]);
  assign t[304] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[305] = (x[66]);
  assign t[306] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[307] = (x[74]);
  assign t[308] = (x[25]);
  assign t[309] = (x[44]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[41]);
  assign t[311] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[312] = (x[85]);
  assign t[313] = (x[52]);
  assign t[314] = (x[49]);
  assign t[315] = (x[33]);
  assign t[316] = (x[62]);
  assign t[317] = (x[59]);
  assign t[318] = (x[68]);
  assign t[319] = (x[65]);
  assign t[31] = t[47] | t[107];
  assign t[320] = (x[76]);
  assign t[321] = (x[73]);
  assign t[322] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[323] = (x[100]);
  assign t[324] = (x[43]);
  assign t[325] = (x[87]);
  assign t[326] = (x[84]);
  assign t[327] = (x[51]);
  assign t[328] = (x[61]);
  assign t[329] = (x[67]);
  assign t[32] = t[105] ? x[30] : x[29];
  assign t[330] = (x[75]);
  assign t[331] = (x[102]);
  assign t[332] = (x[99]);
  assign t[333] = (x[86]);
  assign t[334] = (x[101]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = t[50] ^ t[51];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[35];
  assign t[37] = ~(t[55] & t[56]);
  assign t[38] = t[57] | t[108];
  assign t[39] = t[58] ? x[38] : x[37];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[41];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[109]);
  assign t[46] = ~(t[110]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[69] & t[70]);
  assign t[49] = t[71] | t[111];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[105] ? x[48] : x[47];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = ~(t[74] & t[75]);
  assign t[53] = t[76] | t[112];
  assign t[54] = t[105] ? x[56] : x[55];
  assign t[55] = ~(t[113]);
  assign t[56] = ~(t[114]);
  assign t[57] = ~(t[77] | t[55]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[78] & t[79]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[80] | t[115];
  assign t[61] = ~(t[81] & t[82]);
  assign t[62] = t[83] | t[116];
  assign t[63] = t[18] ? x[72] : x[71];
  assign t[64] = ~(t[84] & t[85]);
  assign t[65] = t[86] | t[117];
  assign t[66] = t[18] ? x[80] : x[79];
  assign t[67] = ~(t[87] & t[88]);
  assign t[68] = ~(t[118]);
  assign t[69] = ~(t[119]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[120]);
  assign t[71] = ~(t[89] | t[69]);
  assign t[72] = ~(t[90] & t[91]);
  assign t[73] = t[92] | t[121];
  assign t[74] = ~(t[122]);
  assign t[75] = ~(t[123]);
  assign t[76] = ~(t[93] | t[74]);
  assign t[77] = ~(t[124]);
  assign t[78] = ~(t[125]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[94] | t[78]);
  assign t[81] = ~(t[127]);
  assign t[82] = ~(t[128]);
  assign t[83] = ~(t[95] | t[81]);
  assign t[84] = ~(t[129]);
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[96] | t[84]);
  assign t[87] = ~(t[97] & t[98]);
  assign t[88] = t[99] | t[131];
  assign t[89] = ~(t[132]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[100] | t[90]);
  assign t[93] = ~(t[135]);
  assign t[94] = ~(t[136]);
  assign t[95] = ~(t[137]);
  assign t[96] = ~(t[138]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[101] | t[97]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [115:0] x;
 output y;

 wire [343:0] t;
  assign t[0] = t[1] ? t[2] : t[111];
  assign t[100] = ~(t[137] & t[136]);
  assign t[101] = ~(t[146]);
  assign t[102] = ~(t[139] & t[138]);
  assign t[103] = ~(t[147]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[109] & t[110]);
  assign t[107] = ~(t[143] & t[142]);
  assign t[108] = ~(t[150]);
  assign t[109] = ~(t[149] & t[148]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = t[193] ^ x[5];
  assign t[153] = t[194] ^ x[13];
  assign t[154] = t[195] ^ x[16];
  assign t[155] = t[196] ^ x[19];
  assign t[156] = t[197] ^ x[22];
  assign t[157] = t[198] ^ x[28];
  assign t[158] = t[199] ^ x[36];
  assign t[159] = t[200] ^ x[39];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[40];
  assign t[161] = t[202] ^ x[46];
  assign t[162] = t[203] ^ x[54];
  assign t[163] = t[204] ^ x[57];
  assign t[164] = t[205] ^ x[58];
  assign t[165] = t[206] ^ x[64];
  assign t[166] = t[207] ^ x[70];
  assign t[167] = t[208] ^ x[78];
  assign t[168] = t[209] ^ x[81];
  assign t[169] = t[210] ^ x[82];
  assign t[16] = ~(t[112] & t[113]);
  assign t[170] = t[211] ^ x[83];
  assign t[171] = t[212] ^ x[89];
  assign t[172] = t[213] ^ x[90];
  assign t[173] = t[214] ^ x[91];
  assign t[174] = t[215] ^ x[92];
  assign t[175] = t[216] ^ x[93];
  assign t[176] = t[217] ^ x[94];
  assign t[177] = t[218] ^ x[95];
  assign t[178] = t[219] ^ x[96];
  assign t[179] = t[220] ^ x[97];
  assign t[17] = ~(t[114] & t[115]);
  assign t[180] = t[221] ^ x[98];
  assign t[181] = t[222] ^ x[104];
  assign t[182] = t[223] ^ x[105];
  assign t[183] = t[224] ^ x[106];
  assign t[184] = t[225] ^ x[107];
  assign t[185] = t[226] ^ x[108];
  assign t[186] = t[227] ^ x[109];
  assign t[187] = t[228] ^ x[110];
  assign t[188] = t[229] ^ x[111];
  assign t[189] = t[230] ^ x[112];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[113];
  assign t[191] = t[232] ^ x[114];
  assign t[192] = t[233] ^ x[115];
  assign t[193] = (~t[234] & t[235]);
  assign t[194] = (~t[236] & t[237]);
  assign t[195] = (~t[238] & t[239]);
  assign t[196] = (~t[240] & t[241]);
  assign t[197] = (~t[242] & t[243]);
  assign t[198] = (~t[244] & t[245]);
  assign t[199] = (~t[246] & t[247]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[244] & t[248]);
  assign t[201] = (~t[244] & t[249]);
  assign t[202] = (~t[250] & t[251]);
  assign t[203] = (~t[252] & t[253]);
  assign t[204] = (~t[246] & t[254]);
  assign t[205] = (~t[246] & t[255]);
  assign t[206] = (~t[256] & t[257]);
  assign t[207] = (~t[258] & t[259]);
  assign t[208] = (~t[260] & t[261]);
  assign t[209] = (~t[244] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[250] & t[263]);
  assign t[211] = (~t[250] & t[264]);
  assign t[212] = (~t[265] & t[266]);
  assign t[213] = (~t[252] & t[267]);
  assign t[214] = (~t[252] & t[268]);
  assign t[215] = (~t[246] & t[269]);
  assign t[216] = (~t[256] & t[270]);
  assign t[217] = (~t[256] & t[271]);
  assign t[218] = (~t[258] & t[272]);
  assign t[219] = (~t[258] & t[273]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[260] & t[274]);
  assign t[221] = (~t[260] & t[275]);
  assign t[222] = (~t[276] & t[277]);
  assign t[223] = (~t[250] & t[278]);
  assign t[224] = (~t[265] & t[279]);
  assign t[225] = (~t[265] & t[280]);
  assign t[226] = (~t[252] & t[281]);
  assign t[227] = (~t[256] & t[282]);
  assign t[228] = (~t[258] & t[283]);
  assign t[229] = (~t[260] & t[284]);
  assign t[22] = t[32] ^ t[26];
  assign t[230] = (~t[276] & t[285]);
  assign t[231] = (~t[276] & t[286]);
  assign t[232] = (~t[265] & t[287]);
  assign t[233] = (~t[276] & t[288]);
  assign t[234] = t[289] ^ x[4];
  assign t[235] = t[290] ^ x[5];
  assign t[236] = t[291] ^ x[12];
  assign t[237] = t[292] ^ x[13];
  assign t[238] = t[293] ^ x[15];
  assign t[239] = t[294] ^ x[16];
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = t[295] ^ x[18];
  assign t[241] = t[296] ^ x[19];
  assign t[242] = t[297] ^ x[21];
  assign t[243] = t[298] ^ x[22];
  assign t[244] = t[299] ^ x[27];
  assign t[245] = t[300] ^ x[28];
  assign t[246] = t[301] ^ x[35];
  assign t[247] = t[302] ^ x[36];
  assign t[248] = t[303] ^ x[39];
  assign t[249] = t[304] ^ x[40];
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = t[305] ^ x[45];
  assign t[251] = t[306] ^ x[46];
  assign t[252] = t[307] ^ x[53];
  assign t[253] = t[308] ^ x[54];
  assign t[254] = t[309] ^ x[57];
  assign t[255] = t[310] ^ x[58];
  assign t[256] = t[311] ^ x[63];
  assign t[257] = t[312] ^ x[64];
  assign t[258] = t[313] ^ x[69];
  assign t[259] = t[314] ^ x[70];
  assign t[25] = ~(t[114]);
  assign t[260] = t[315] ^ x[77];
  assign t[261] = t[316] ^ x[78];
  assign t[262] = t[317] ^ x[81];
  assign t[263] = t[318] ^ x[82];
  assign t[264] = t[319] ^ x[83];
  assign t[265] = t[320] ^ x[88];
  assign t[266] = t[321] ^ x[89];
  assign t[267] = t[322] ^ x[90];
  assign t[268] = t[323] ^ x[91];
  assign t[269] = t[324] ^ x[92];
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = t[325] ^ x[93];
  assign t[271] = t[326] ^ x[94];
  assign t[272] = t[327] ^ x[95];
  assign t[273] = t[328] ^ x[96];
  assign t[274] = t[329] ^ x[97];
  assign t[275] = t[330] ^ x[98];
  assign t[276] = t[331] ^ x[103];
  assign t[277] = t[332] ^ x[104];
  assign t[278] = t[333] ^ x[105];
  assign t[279] = t[334] ^ x[106];
  assign t[27] = t[39] ^ t[40];
  assign t[280] = t[335] ^ x[107];
  assign t[281] = t[336] ^ x[108];
  assign t[282] = t[337] ^ x[109];
  assign t[283] = t[338] ^ x[110];
  assign t[284] = t[339] ^ x[111];
  assign t[285] = t[340] ^ x[112];
  assign t[286] = t[341] ^ x[113];
  assign t[287] = t[342] ^ x[114];
  assign t[288] = t[343] ^ x[115];
  assign t[289] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[290] = (x[2]);
  assign t[291] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[292] = (x[11]);
  assign t[293] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[294] = (x[14]);
  assign t[295] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[296] = (x[17]);
  assign t[297] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[298] = (x[20]);
  assign t[299] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[24]);
  assign t[301] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[302] = (x[32]);
  assign t[303] = (x[26]);
  assign t[304] = (x[23]);
  assign t[305] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[306] = (x[42]);
  assign t[307] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[308] = (x[50]);
  assign t[309] = (x[34]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[31]);
  assign t[311] = (x[59] & ~x[60] & ~x[61] & ~x[62]) | (~x[59] & x[60] & ~x[61] & ~x[62]) | (~x[59] & ~x[60] & x[61] & ~x[62]) | (~x[59] & ~x[60] & ~x[61] & x[62]) | (x[59] & x[60] & x[61] & ~x[62]) | (x[59] & x[60] & ~x[61] & x[62]) | (x[59] & ~x[60] & x[61] & x[62]) | (~x[59] & x[60] & x[61] & x[62]);
  assign t[312] = (x[60]);
  assign t[313] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[314] = (x[66]);
  assign t[315] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[316] = (x[74]);
  assign t[317] = (x[25]);
  assign t[318] = (x[44]);
  assign t[319] = (x[41]);
  assign t[31] = ~(t[47] & t[116]);
  assign t[320] = (x[84] & ~x[85] & ~x[86] & ~x[87]) | (~x[84] & x[85] & ~x[86] & ~x[87]) | (~x[84] & ~x[85] & x[86] & ~x[87]) | (~x[84] & ~x[85] & ~x[86] & x[87]) | (x[84] & x[85] & x[86] & ~x[87]) | (x[84] & x[85] & ~x[86] & x[87]) | (x[84] & ~x[85] & x[86] & x[87]) | (~x[84] & x[85] & x[86] & x[87]);
  assign t[321] = (x[85]);
  assign t[322] = (x[52]);
  assign t[323] = (x[49]);
  assign t[324] = (x[33]);
  assign t[325] = (x[62]);
  assign t[326] = (x[59]);
  assign t[327] = (x[68]);
  assign t[328] = (x[65]);
  assign t[329] = (x[76]);
  assign t[32] = t[114] ? x[30] : x[29];
  assign t[330] = (x[73]);
  assign t[331] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[332] = (x[100]);
  assign t[333] = (x[43]);
  assign t[334] = (x[87]);
  assign t[335] = (x[84]);
  assign t[336] = (x[51]);
  assign t[337] = (x[61]);
  assign t[338] = (x[67]);
  assign t[339] = (x[75]);
  assign t[33] = ~(t[48] & t[49]);
  assign t[340] = (x[102]);
  assign t[341] = (x[99]);
  assign t[342] = (x[86]);
  assign t[343] = (x[101]);
  assign t[34] = t[50] ^ t[51];
  assign t[35] = ~(t[52] & t[53]);
  assign t[36] = t[54] ^ t[35];
  assign t[37] = ~(t[55] & t[56]);
  assign t[38] = ~(t[57] & t[117]);
  assign t[39] = t[58] ? x[38] : x[37];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[59] & t[60]);
  assign t[41] = ~(t[61] & t[62]);
  assign t[42] = t[63] ^ t[41];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[118]);
  assign t[46] = ~(t[119]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = ~(t[70] & t[71]);
  assign t[49] = ~(t[72] & t[120]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[114] ? x[48] : x[47];
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[76]);
  assign t[53] = ~(t[77] & t[121]);
  assign t[54] = t[114] ? x[56] : x[55];
  assign t[55] = ~(t[122]);
  assign t[56] = ~(t[123]);
  assign t[57] = ~(t[78] & t[79]);
  assign t[58] = ~(t[25]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[82] & t[124]);
  assign t[61] = ~(t[83] & t[84]);
  assign t[62] = ~(t[85] & t[125]);
  assign t[63] = t[18] ? x[72] : x[71];
  assign t[64] = ~(t[86] & t[87]);
  assign t[65] = ~(t[88] & t[126]);
  assign t[66] = t[18] ? x[80] : x[79];
  assign t[67] = ~(t[89] & t[90]);
  assign t[68] = ~(t[119] & t[118]);
  assign t[69] = ~(t[127]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[128]);
  assign t[71] = ~(t[129]);
  assign t[72] = ~(t[91] & t[92]);
  assign t[73] = ~(t[93] & t[94]);
  assign t[74] = ~(t[95] & t[130]);
  assign t[75] = ~(t[131]);
  assign t[76] = ~(t[132]);
  assign t[77] = ~(t[96] & t[97]);
  assign t[78] = ~(t[123] & t[122]);
  assign t[79] = ~(t[133]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[134]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[98] & t[99]);
  assign t[83] = ~(t[136]);
  assign t[84] = ~(t[137]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[102] & t[103]);
  assign t[89] = ~(t[104] & t[105]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[106] & t[140]);
  assign t[91] = ~(t[129] & t[128]);
  assign t[92] = ~(t[141]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[143]);
  assign t[95] = ~(t[107] & t[108]);
  assign t[96] = ~(t[132] & t[131]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[135] & t[134]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [106:0] x;
 output y;

 wire [280:0] t;
  assign t[0] = t[1] ? t[2] : t[93];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = t[157] ^ x[5];
  assign t[126] = t[158] ^ x[13];
  assign t[127] = t[159] ^ x[16];
  assign t[128] = t[160] ^ x[19];
  assign t[129] = t[161] ^ x[22];
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = t[162] ^ x[28];
  assign t[131] = t[163] ^ x[29];
  assign t[132] = t[164] ^ x[37];
  assign t[133] = t[165] ^ x[38];
  assign t[134] = t[166] ^ x[41];
  assign t[135] = t[167] ^ x[47];
  assign t[136] = t[168] ^ x[48];
  assign t[137] = t[169] ^ x[56];
  assign t[138] = t[170] ^ x[57];
  assign t[139] = t[171] ^ x[60];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[66];
  assign t[141] = t[173] ^ x[67];
  assign t[142] = t[174] ^ x[73];
  assign t[143] = t[175] ^ x[74];
  assign t[144] = t[176] ^ x[82];
  assign t[145] = t[177] ^ x[83];
  assign t[146] = t[178] ^ x[86];
  assign t[147] = t[179] ^ x[87];
  assign t[148] = t[180] ^ x[93];
  assign t[149] = t[181] ^ x[94];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[95];
  assign t[151] = t[183] ^ x[96];
  assign t[152] = t[184] ^ x[102];
  assign t[153] = t[185] ^ x[103];
  assign t[154] = t[186] ^ x[104];
  assign t[155] = t[187] ^ x[105];
  assign t[156] = t[188] ^ x[106];
  assign t[157] = (~t[189] & t[190]);
  assign t[158] = (~t[191] & t[192]);
  assign t[159] = (~t[193] & t[194]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (~t[195] & t[196]);
  assign t[161] = (~t[197] & t[198]);
  assign t[162] = (~t[199] & t[200]);
  assign t[163] = (~t[199] & t[201]);
  assign t[164] = (~t[202] & t[203]);
  assign t[165] = (~t[202] & t[204]);
  assign t[166] = (~t[199] & t[205]);
  assign t[167] = (~t[206] & t[207]);
  assign t[168] = (~t[206] & t[208]);
  assign t[169] = (~t[209] & t[210]);
  assign t[16] = ~(t[94] & t[95]);
  assign t[170] = (~t[209] & t[211]);
  assign t[171] = (~t[202] & t[212]);
  assign t[172] = (~t[213] & t[214]);
  assign t[173] = (~t[213] & t[215]);
  assign t[174] = (~t[216] & t[217]);
  assign t[175] = (~t[216] & t[218]);
  assign t[176] = (~t[219] & t[220]);
  assign t[177] = (~t[219] & t[221]);
  assign t[178] = (~t[206] & t[222]);
  assign t[179] = (~t[209] & t[223]);
  assign t[17] = ~(t[96] & t[97]);
  assign t[180] = (~t[224] & t[225]);
  assign t[181] = (~t[224] & t[226]);
  assign t[182] = (~t[213] & t[227]);
  assign t[183] = (~t[216] & t[228]);
  assign t[184] = (~t[229] & t[230]);
  assign t[185] = (~t[229] & t[231]);
  assign t[186] = (~t[219] & t[232]);
  assign t[187] = (~t[224] & t[233]);
  assign t[188] = (~t[229] & t[234]);
  assign t[189] = t[235] ^ x[4];
  assign t[18] = ~(t[25]);
  assign t[190] = t[236] ^ x[5];
  assign t[191] = t[237] ^ x[12];
  assign t[192] = t[238] ^ x[13];
  assign t[193] = t[239] ^ x[15];
  assign t[194] = t[240] ^ x[16];
  assign t[195] = t[241] ^ x[18];
  assign t[196] = t[242] ^ x[19];
  assign t[197] = t[243] ^ x[21];
  assign t[198] = t[244] ^ x[22];
  assign t[199] = t[245] ^ x[27];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[246] ^ x[28];
  assign t[201] = t[247] ^ x[29];
  assign t[202] = t[248] ^ x[36];
  assign t[203] = t[249] ^ x[37];
  assign t[204] = t[250] ^ x[38];
  assign t[205] = t[251] ^ x[41];
  assign t[206] = t[252] ^ x[46];
  assign t[207] = t[253] ^ x[47];
  assign t[208] = t[254] ^ x[48];
  assign t[209] = t[255] ^ x[55];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[256] ^ x[56];
  assign t[211] = t[257] ^ x[57];
  assign t[212] = t[258] ^ x[60];
  assign t[213] = t[259] ^ x[65];
  assign t[214] = t[260] ^ x[66];
  assign t[215] = t[261] ^ x[67];
  assign t[216] = t[262] ^ x[72];
  assign t[217] = t[263] ^ x[73];
  assign t[218] = t[264] ^ x[74];
  assign t[219] = t[265] ^ x[81];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[266] ^ x[82];
  assign t[221] = t[267] ^ x[83];
  assign t[222] = t[268] ^ x[86];
  assign t[223] = t[269] ^ x[87];
  assign t[224] = t[270] ^ x[92];
  assign t[225] = t[271] ^ x[93];
  assign t[226] = t[272] ^ x[94];
  assign t[227] = t[273] ^ x[95];
  assign t[228] = t[274] ^ x[96];
  assign t[229] = t[275] ^ x[101];
  assign t[22] = t[32] ^ t[26];
  assign t[230] = t[276] ^ x[102];
  assign t[231] = t[277] ^ x[103];
  assign t[232] = t[278] ^ x[104];
  assign t[233] = t[279] ^ x[105];
  assign t[234] = t[280] ^ x[106];
  assign t[235] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[236] = (x[1]);
  assign t[237] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[238] = (x[11]);
  assign t[239] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[23] = x[7] ? t[34] : t[33];
  assign t[240] = (x[14]);
  assign t[241] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[242] = (x[17]);
  assign t[243] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[244] = (x[20]);
  assign t[245] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[246] = (x[25]);
  assign t[247] = (x[23]);
  assign t[248] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[249] = (x[34]);
  assign t[24] = x[7] ? t[36] : t[35];
  assign t[250] = (x[32]);
  assign t[251] = (x[26]);
  assign t[252] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[253] = (x[44]);
  assign t[254] = (x[42]);
  assign t[255] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[256] = (x[53]);
  assign t[257] = (x[51]);
  assign t[258] = (x[35]);
  assign t[259] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[25] = ~(t[96]);
  assign t[260] = (x[63]);
  assign t[261] = (x[61]);
  assign t[262] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[263] = (x[70]);
  assign t[264] = (x[68]);
  assign t[265] = (x[77] & ~x[78] & ~x[79] & ~x[80]) | (~x[77] & x[78] & ~x[79] & ~x[80]) | (~x[77] & ~x[78] & x[79] & ~x[80]) | (~x[77] & ~x[78] & ~x[79] & x[80]) | (x[77] & x[78] & x[79] & ~x[80]) | (x[77] & x[78] & ~x[79] & x[80]) | (x[77] & ~x[78] & x[79] & x[80]) | (~x[77] & x[78] & x[79] & x[80]);
  assign t[266] = (x[79]);
  assign t[267] = (x[77]);
  assign t[268] = (x[45]);
  assign t[269] = (x[54]);
  assign t[26] = ~(t[37] & t[38]);
  assign t[270] = (x[88] & ~x[89] & ~x[90] & ~x[91]) | (~x[88] & x[89] & ~x[90] & ~x[91]) | (~x[88] & ~x[89] & x[90] & ~x[91]) | (~x[88] & ~x[89] & ~x[90] & x[91]) | (x[88] & x[89] & x[90] & ~x[91]) | (x[88] & x[89] & ~x[90] & x[91]) | (x[88] & ~x[89] & x[90] & x[91]) | (~x[88] & x[89] & x[90] & x[91]);
  assign t[271] = (x[90]);
  assign t[272] = (x[88]);
  assign t[273] = (x[64]);
  assign t[274] = (x[71]);
  assign t[275] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[276] = (x[99]);
  assign t[277] = (x[97]);
  assign t[278] = (x[80]);
  assign t[279] = (x[91]);
  assign t[27] = t[39] ^ t[40];
  assign t[280] = (x[100]);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[98] & t[45]);
  assign t[31] = ~(t[99] & t[46]);
  assign t[32] = t[96] ? x[31] : x[30];
  assign t[33] = ~(t[47] & t[48]);
  assign t[34] = t[49] ^ t[33];
  assign t[35] = ~(t[50] & t[51]);
  assign t[36] = t[52] ^ t[53];
  assign t[37] = ~(t[100] & t[54]);
  assign t[38] = ~(t[101] & t[55]);
  assign t[39] = t[56] ? x[40] : x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[57] & t[58]);
  assign t[41] = ~(t[59] & t[60]);
  assign t[42] = t[61] ^ t[62];
  assign t[43] = ~(t[63] & t[64]);
  assign t[44] = t[65] ^ t[43];
  assign t[45] = ~(t[102]);
  assign t[46] = ~(t[102] & t[66]);
  assign t[47] = ~(t[103] & t[67]);
  assign t[48] = ~(t[104] & t[68]);
  assign t[49] = t[96] ? x[50] : x[49];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[105] & t[69]);
  assign t[51] = ~(t[106] & t[70]);
  assign t[52] = t[96] ? x[59] : x[58];
  assign t[53] = ~(t[71] & t[72]);
  assign t[54] = ~(t[107]);
  assign t[55] = ~(t[107] & t[73]);
  assign t[56] = ~(t[25]);
  assign t[57] = ~(t[108] & t[74]);
  assign t[58] = ~(t[109] & t[75]);
  assign t[59] = ~(t[110] & t[76]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[111] & t[77]);
  assign t[61] = t[18] ? x[76] : x[75];
  assign t[62] = ~(t[78] & t[79]);
  assign t[63] = ~(t[112] & t[80]);
  assign t[64] = ~(t[113] & t[81]);
  assign t[65] = t[18] ? x[85] : x[84];
  assign t[66] = ~(t[98]);
  assign t[67] = ~(t[114]);
  assign t[68] = ~(t[114] & t[82]);
  assign t[69] = ~(t[115]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[115] & t[83]);
  assign t[71] = ~(t[116] & t[84]);
  assign t[72] = ~(t[117] & t[85]);
  assign t[73] = ~(t[100]);
  assign t[74] = ~(t[118]);
  assign t[75] = ~(t[118] & t[86]);
  assign t[76] = ~(t[119]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121] & t[89]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[122]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[103]);
  assign t[83] = ~(t[105]);
  assign t[84] = ~(t[123]);
  assign t[85] = ~(t[123] & t[91]);
  assign t[86] = ~(t[108]);
  assign t[87] = ~(t[110]);
  assign t[88] = ~(t[124]);
  assign t[89] = ~(t[124] & t[92]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[112]);
  assign t[91] = ~(t[116]);
  assign t[92] = ~(t[120]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [115:0] x;
 output y;

 wire [433:0] t;
  assign t[0] = t[1] ? t[2] : t[201];
  assign t[100] = ~(t[223]);
  assign t[101] = ~(t[212] | t[213]);
  assign t[102] = ~(t[224]);
  assign t[103] = ~(t[225]);
  assign t[104] = ~(t[140] | t[141]);
  assign t[105] = ~(t[48]);
  assign t[106] = ~(t[129] | t[142]);
  assign t[107] = ~(t[127]);
  assign t[108] = ~(t[226]);
  assign t[109] = ~(t[227]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[143] | t[144]);
  assign t[111] = t[30] ? x[94] : x[93];
  assign t[112] = ~(t[145] & t[146]);
  assign t[113] = ~(t[228]);
  assign t[114] = ~(t[229]);
  assign t[115] = ~(t[147] | t[148]);
  assign t[116] = ~(t[149] | t[150]);
  assign t[117] = ~(t[230] | t[151]);
  assign t[118] = t[30] ? x[104] : x[103];
  assign t[119] = ~(t[83] & t[152]);
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[204]);
  assign t[121] = ~(t[205] & t[153]);
  assign t[122] = ~(x[7] & t[154]);
  assign t[123] = ~(t[155] & t[205]);
  assign t[124] = ~(t[156] & t[157]);
  assign t[125] = ~(t[120] | t[158]);
  assign t[126] = ~(t[120] | t[159]);
  assign t[127] = ~(t[79] | t[160]);
  assign t[128] = ~(t[161] & t[162]);
  assign t[129] = ~(t[79] | t[163]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = ~(t[231]);
  assign t[131] = ~(t[218] | t[219]);
  assign t[132] = ~(t[232]);
  assign t[133] = ~(t[233]);
  assign t[134] = ~(t[164] | t[165]);
  assign t[135] = ~(t[138] | t[166]);
  assign t[136] = ~(t[234]);
  assign t[137] = ~(t[221] | t[222]);
  assign t[138] = ~(t[167] & t[168]);
  assign t[139] = ~(t[169] & t[31]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[235]);
  assign t[141] = ~(t[224] | t[225]);
  assign t[142] = ~(t[170] & t[83]);
  assign t[143] = ~(t[236]);
  assign t[144] = ~(t[226] | t[227]);
  assign t[145] = ~(t[171] | t[126]);
  assign t[146] = ~(t[172] | t[173]);
  assign t[147] = ~(t[237]);
  assign t[148] = ~(t[228] | t[229]);
  assign t[149] = ~(t[238]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[239]);
  assign t[151] = ~(t[174] | t[175]);
  assign t[152] = ~(t[176] | t[177]);
  assign t[153] = ~(x[7] | t[178]);
  assign t[154] = ~(t[203] | t[205]);
  assign t[155] = ~(x[7] | t[203]);
  assign t[156] = x[7] & t[203];
  assign t[157] = ~(t[205]);
  assign t[158] = t[202] ? t[124] : t[179];
  assign t[159] = t[202] ? t[180] : t[122];
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = t[202] ? t[179] : t[181];
  assign t[161] = ~(t[182] | t[49]);
  assign t[162] = ~(t[51] & t[183]);
  assign t[163] = t[202] ? t[184] : t[180];
  assign t[164] = ~(t[240]);
  assign t[165] = ~(t[232] | t[233]);
  assign t[166] = ~(t[185] & t[186]);
  assign t[167] = ~(t[82] & t[187]);
  assign t[168] = ~(t[188] & t[189]);
  assign t[169] = ~(t[127] | t[190]);
  assign t[16] = ~(t[202] & t[203]);
  assign t[170] = ~(t[182] | t[176]);
  assign t[171] = ~(t[120] | t[191]);
  assign t[172] = ~(t[87]);
  assign t[173] = ~(t[79] | t[192]);
  assign t[174] = ~(t[241]);
  assign t[175] = ~(t[238] | t[239]);
  assign t[176] = ~(t[193] & t[194]);
  assign t[177] = ~(t[162] & t[186]);
  assign t[178] = ~(t[203]);
  assign t[179] = ~(t[155] & t[157]);
  assign t[17] = ~(t[204] & t[205]);
  assign t[180] = ~(t[153] & t[157]);
  assign t[181] = ~(t[156] & t[205]);
  assign t[182] = ~(t[79] | t[195]);
  assign t[183] = t[155] | t[156];
  assign t[184] = ~(x[7] & t[188]);
  assign t[185] = ~(t[126]);
  assign t[186] = t[120] | t[196];
  assign t[187] = ~(t[121] & t[184]);
  assign t[188] = ~(t[203] | t[157]);
  assign t[189] = t[79] & t[202];
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = ~(t[79] | t[197]);
  assign t[191] = t[202] ? t[179] : t[124];
  assign t[192] = t[202] ? t[121] : t[122];
  assign t[193] = ~(t[171] | t[198]);
  assign t[194] = ~(t[120] & t[199]);
  assign t[195] = t[202] ? t[181] : t[179];
  assign t[196] = t[202] ? t[122] : t[180];
  assign t[197] = t[202] ? t[123] : t[124];
  assign t[198] = ~(t[79] | t[200]);
  assign t[199] = ~(t[122] & t[121]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[202] ? t[180] : t[184];
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = (t[280]);
  assign t[23] = ~(t[26] ^ t[35]);
  assign t[240] = (t[281]);
  assign t[241] = (t[282]);
  assign t[242] = t[283] ^ x[5];
  assign t[243] = t[284] ^ x[13];
  assign t[244] = t[285] ^ x[16];
  assign t[245] = t[286] ^ x[19];
  assign t[246] = t[287] ^ x[22];
  assign t[247] = t[288] ^ x[28];
  assign t[248] = t[289] ^ x[34];
  assign t[249] = t[290] ^ x[35];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[291] ^ x[36];
  assign t[251] = t[292] ^ x[44];
  assign t[252] = t[293] ^ x[50];
  assign t[253] = t[294] ^ x[51];
  assign t[254] = t[295] ^ x[52];
  assign t[255] = t[296] ^ x[58];
  assign t[256] = t[297] ^ x[66];
  assign t[257] = t[298] ^ x[72];
  assign t[258] = t[299] ^ x[73];
  assign t[259] = t[300] ^ x[74];
  assign t[25] = x[7] ? t[39] : t[38];
  assign t[260] = t[301] ^ x[75];
  assign t[261] = t[302] ^ x[81];
  assign t[262] = t[303] ^ x[84];
  assign t[263] = t[304] ^ x[85];
  assign t[264] = t[305] ^ x[88];
  assign t[265] = t[306] ^ x[89];
  assign t[266] = t[307] ^ x[90];
  assign t[267] = t[308] ^ x[91];
  assign t[268] = t[309] ^ x[92];
  assign t[269] = t[310] ^ x[95];
  assign t[26] = ~(t[40] | t[41]);
  assign t[270] = t[311] ^ x[96];
  assign t[271] = t[312] ^ x[102];
  assign t[272] = t[313] ^ x[105];
  assign t[273] = t[314] ^ x[106];
  assign t[274] = t[315] ^ x[107];
  assign t[275] = t[316] ^ x[108];
  assign t[276] = t[317] ^ x[109];
  assign t[277] = t[318] ^ x[110];
  assign t[278] = t[319] ^ x[111];
  assign t[279] = t[320] ^ x[112];
  assign t[27] = ~(t[42] ^ t[43]);
  assign t[280] = t[321] ^ x[113];
  assign t[281] = t[322] ^ x[114];
  assign t[282] = t[323] ^ x[115];
  assign t[283] = (~t[324] & t[325]);
  assign t[284] = (~t[326] & t[327]);
  assign t[285] = (~t[328] & t[329]);
  assign t[286] = (~t[330] & t[331]);
  assign t[287] = (~t[332] & t[333]);
  assign t[288] = (~t[334] & t[335]);
  assign t[289] = (~t[336] & t[337]);
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = (~t[334] & t[338]);
  assign t[291] = (~t[334] & t[339]);
  assign t[292] = (~t[340] & t[341]);
  assign t[293] = (~t[342] & t[343]);
  assign t[294] = (~t[336] & t[344]);
  assign t[295] = (~t[336] & t[345]);
  assign t[296] = (~t[346] & t[347]);
  assign t[297] = (~t[348] & t[349]);
  assign t[298] = (~t[350] & t[351]);
  assign t[299] = (~t[334] & t[352]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[340] & t[353]);
  assign t[301] = (~t[340] & t[354]);
  assign t[302] = (~t[355] & t[356]);
  assign t[303] = (~t[342] & t[357]);
  assign t[304] = (~t[342] & t[358]);
  assign t[305] = (~t[336] & t[359]);
  assign t[306] = (~t[346] & t[360]);
  assign t[307] = (~t[346] & t[361]);
  assign t[308] = (~t[348] & t[362]);
  assign t[309] = (~t[348] & t[363]);
  assign t[30] = ~(t[48]);
  assign t[310] = (~t[350] & t[364]);
  assign t[311] = (~t[350] & t[365]);
  assign t[312] = (~t[366] & t[367]);
  assign t[313] = (~t[340] & t[368]);
  assign t[314] = (~t[355] & t[369]);
  assign t[315] = (~t[355] & t[370]);
  assign t[316] = (~t[342] & t[371]);
  assign t[317] = (~t[346] & t[372]);
  assign t[318] = (~t[348] & t[373]);
  assign t[319] = (~t[350] & t[374]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (~t[366] & t[375]);
  assign t[321] = (~t[366] & t[376]);
  assign t[322] = (~t[355] & t[377]);
  assign t[323] = (~t[366] & t[378]);
  assign t[324] = t[379] ^ x[4];
  assign t[325] = t[380] ^ x[5];
  assign t[326] = t[381] ^ x[12];
  assign t[327] = t[382] ^ x[13];
  assign t[328] = t[383] ^ x[15];
  assign t[329] = t[384] ^ x[16];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[385] ^ x[18];
  assign t[331] = t[386] ^ x[19];
  assign t[332] = t[387] ^ x[21];
  assign t[333] = t[388] ^ x[22];
  assign t[334] = t[389] ^ x[27];
  assign t[335] = t[390] ^ x[28];
  assign t[336] = t[391] ^ x[33];
  assign t[337] = t[392] ^ x[34];
  assign t[338] = t[393] ^ x[35];
  assign t[339] = t[394] ^ x[36];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[395] ^ x[43];
  assign t[341] = t[396] ^ x[44];
  assign t[342] = t[397] ^ x[49];
  assign t[343] = t[398] ^ x[50];
  assign t[344] = t[399] ^ x[51];
  assign t[345] = t[400] ^ x[52];
  assign t[346] = t[401] ^ x[57];
  assign t[347] = t[402] ^ x[58];
  assign t[348] = t[403] ^ x[65];
  assign t[349] = t[404] ^ x[66];
  assign t[34] = ~(t[206] | t[55]);
  assign t[350] = t[405] ^ x[71];
  assign t[351] = t[406] ^ x[72];
  assign t[352] = t[407] ^ x[73];
  assign t[353] = t[408] ^ x[74];
  assign t[354] = t[409] ^ x[75];
  assign t[355] = t[410] ^ x[80];
  assign t[356] = t[411] ^ x[81];
  assign t[357] = t[412] ^ x[84];
  assign t[358] = t[413] ^ x[85];
  assign t[359] = t[414] ^ x[88];
  assign t[35] = ~(t[56] ^ t[57]);
  assign t[360] = t[415] ^ x[89];
  assign t[361] = t[416] ^ x[90];
  assign t[362] = t[417] ^ x[91];
  assign t[363] = t[418] ^ x[92];
  assign t[364] = t[419] ^ x[95];
  assign t[365] = t[420] ^ x[96];
  assign t[366] = t[421] ^ x[101];
  assign t[367] = t[422] ^ x[102];
  assign t[368] = t[423] ^ x[105];
  assign t[369] = t[424] ^ x[106];
  assign t[36] = ~(t[58] | t[59]);
  assign t[370] = t[425] ^ x[107];
  assign t[371] = t[426] ^ x[108];
  assign t[372] = t[427] ^ x[109];
  assign t[373] = t[428] ^ x[110];
  assign t[374] = t[429] ^ x[111];
  assign t[375] = t[430] ^ x[112];
  assign t[376] = t[431] ^ x[113];
  assign t[377] = t[432] ^ x[114];
  assign t[378] = t[433] ^ x[115];
  assign t[379] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = ~(t[60] ^ t[61]);
  assign t[380] = (x[0]);
  assign t[381] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[382] = (x[11]);
  assign t[383] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[384] = (x[14]);
  assign t[385] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[386] = (x[17]);
  assign t[387] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[388] = (x[20]);
  assign t[389] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[38] = ~(t[62] | t[63]);
  assign t[390] = (x[24]);
  assign t[391] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[392] = (x[30]);
  assign t[393] = (x[25]);
  assign t[394] = (x[26]);
  assign t[395] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[396] = (x[40]);
  assign t[397] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[398] = (x[46]);
  assign t[399] = (x[31]);
  assign t[39] = ~(t[38] ^ t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[32]);
  assign t[401] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[402] = (x[54]);
  assign t[403] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[404] = (x[62]);
  assign t[405] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[406] = (x[68]);
  assign t[407] = (x[23]);
  assign t[408] = (x[41]);
  assign t[409] = (x[42]);
  assign t[40] = ~(t[65] | t[66]);
  assign t[410] = (x[76] & ~x[77] & ~x[78] & ~x[79]) | (~x[76] & x[77] & ~x[78] & ~x[79]) | (~x[76] & ~x[77] & x[78] & ~x[79]) | (~x[76] & ~x[77] & ~x[78] & x[79]) | (x[76] & x[77] & x[78] & ~x[79]) | (x[76] & x[77] & ~x[78] & x[79]) | (x[76] & ~x[77] & x[78] & x[79]) | (~x[76] & x[77] & x[78] & x[79]);
  assign t[411] = (x[77]);
  assign t[412] = (x[47]);
  assign t[413] = (x[48]);
  assign t[414] = (x[29]);
  assign t[415] = (x[55]);
  assign t[416] = (x[56]);
  assign t[417] = (x[63]);
  assign t[418] = (x[64]);
  assign t[419] = (x[69]);
  assign t[41] = ~(t[207] | t[67]);
  assign t[420] = (x[70]);
  assign t[421] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[422] = (x[98]);
  assign t[423] = (x[39]);
  assign t[424] = (x[78]);
  assign t[425] = (x[79]);
  assign t[426] = (x[45]);
  assign t[427] = (x[53]);
  assign t[428] = (x[61]);
  assign t[429] = (x[67]);
  assign t[42] = ~(t[68] | t[69]);
  assign t[430] = (x[99]);
  assign t[431] = (x[100]);
  assign t[432] = (x[76]);
  assign t[433] = (x[97]);
  assign t[43] = ~(t[70] ^ t[71]);
  assign t[44] = ~(t[72] | t[73]);
  assign t[45] = ~(t[44] ^ t[74]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[48] = ~(t[204]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[79] | t[81]);
  assign t[51] = t[205] & t[82];
  assign t[52] = ~(t[83]);
  assign t[53] = ~(t[208]);
  assign t[54] = ~(t[209]);
  assign t[55] = ~(t[84] | t[85]);
  assign t[56] = t[204] ? x[38] : x[37];
  assign t[57] = ~(t[86] & t[87]);
  assign t[58] = ~(t[88] | t[89]);
  assign t[59] = ~(t[210] | t[90]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[91] | t[92]);
  assign t[61] = ~(t[93] ^ t[94]);
  assign t[62] = ~(t[95] | t[96]);
  assign t[63] = ~(t[211] | t[97]);
  assign t[64] = ~(t[98] ^ t[99]);
  assign t[65] = ~(t[212]);
  assign t[66] = ~(t[213]);
  assign t[67] = ~(t[100] | t[101]);
  assign t[68] = ~(t[102] | t[103]);
  assign t[69] = ~(t[214] | t[104]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[105] ? x[60] : x[59];
  assign t[71] = ~(t[106] & t[107]);
  assign t[72] = ~(t[108] | t[109]);
  assign t[73] = ~(t[215] | t[110]);
  assign t[74] = ~(t[111] ^ t[112]);
  assign t[75] = ~(t[113] | t[114]);
  assign t[76] = ~(t[216] | t[115]);
  assign t[77] = ~(t[116] | t[117]);
  assign t[78] = ~(t[118] ^ t[119]);
  assign t[79] = ~(t[120]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[202] ? t[122] : t[121];
  assign t[81] = t[202] ? t[124] : t[123];
  assign t[82] = ~(t[120] | t[202]);
  assign t[83] = ~(t[125] | t[126]);
  assign t[84] = ~(t[217]);
  assign t[85] = ~(t[208] | t[209]);
  assign t[86] = ~(t[127] | t[128]);
  assign t[87] = ~(t[129] | t[50]);
  assign t[88] = ~(t[218]);
  assign t[89] = ~(t[219]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[130] | t[131]);
  assign t[91] = ~(t[132] | t[133]);
  assign t[92] = ~(t[220] | t[134]);
  assign t[93] = t[105] ? x[83] : x[82];
  assign t[94] = ~(t[135] & t[107]);
  assign t[95] = ~(t[221]);
  assign t[96] = ~(t[222]);
  assign t[97] = ~(t[136] | t[137]);
  assign t[98] = t[204] ? x[87] : x[86];
  assign t[99] = t[138] | t[139];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [163:0] x;
 output y;

 wire [631:0] t;
  assign t[0] = t[1] ? t[2] : t[384];
  assign t[100] = ~(t[140] | t[141]);
  assign t[101] = t[137] ? x[83] : x[82];
  assign t[102] = ~(t[142] & t[106]);
  assign t[103] = ~(t[407]);
  assign t[104] = ~(t[396] | t[397]);
  assign t[105] = ~(t[125] | t[50]);
  assign t[106] = ~(t[143] | t[139]);
  assign t[107] = ~(t[408]);
  assign t[108] = ~(t[409]);
  assign t[109] = ~(t[144] | t[145]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[146] | t[147]);
  assign t[111] = ~(t[410] | t[148]);
  assign t[112] = t[30] ? x[94] : x[93];
  assign t[113] = ~(t[149] & t[150]);
  assign t[114] = ~(t[411]);
  assign t[115] = ~(t[412]);
  assign t[116] = ~(t[151] | t[152]);
  assign t[117] = ~(t[153] | t[154]);
  assign t[118] = ~(t[413] | t[155]);
  assign t[119] = t[137] ? x[104] : x[103];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[156] & t[157]);
  assign t[121] = ~(t[158] & t[159]);
  assign t[122] = ~(t[160] & t[159]);
  assign t[123] = ~(x[7] & t[161]);
  assign t[124] = ~(t[162] & t[159]);
  assign t[125] = ~(t[79] | t[163]);
  assign t[126] = ~(t[164] | t[165]);
  assign t[127] = ~(t[123] & t[166]);
  assign t[128] = t[388] & t[167];
  assign t[129] = t[158] | t[160];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[385] ? t[123] : t[124];
  assign t[131] = ~(t[414]);
  assign t[132] = ~(t[401] | t[402]);
  assign t[133] = ~(t[168] & t[169]);
  assign t[134] = t[139] | t[170];
  assign t[135] = ~(t[415]);
  assign t[136] = ~(t[403] | t[404]);
  assign t[137] = ~(t[48]);
  assign t[138] = ~(t[31] & t[169]);
  assign t[139] = ~(t[164] | t[171]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[416]);
  assign t[141] = ~(t[405] | t[406]);
  assign t[142] = ~(t[172]);
  assign t[143] = ~(t[173]);
  assign t[144] = ~(t[417]);
  assign t[145] = ~(t[408] | t[409]);
  assign t[146] = ~(t[418]);
  assign t[147] = ~(t[419]);
  assign t[148] = ~(t[174] | t[175]);
  assign t[149] = ~(t[176] | t[177]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[128] | t[178]);
  assign t[151] = ~(t[420]);
  assign t[152] = ~(t[411] | t[412]);
  assign t[153] = ~(t[421]);
  assign t[154] = ~(t[422]);
  assign t[155] = ~(t[179] | t[180]);
  assign t[156] = ~(t[181] | t[182]);
  assign t[157] = ~(t[183]);
  assign t[158] = ~(x[7] | t[386]);
  assign t[159] = ~(t[388]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = x[7] & t[386];
  assign t[161] = ~(t[386] | t[388]);
  assign t[162] = ~(x[7] | t[184]);
  assign t[163] = t[385] ? t[121] : t[122];
  assign t[164] = ~(t[79]);
  assign t[165] = t[385] ? t[124] : t[185];
  assign t[166] = ~(t[388] & t[162]);
  assign t[167] = ~(t[79] | t[385]);
  assign t[168] = ~(t[167] & t[186]);
  assign t[169] = ~(t[187] & t[188]);
  assign t[16] = ~(t[385] & t[386]);
  assign t[170] = ~(t[164] | t[189]);
  assign t[171] = t[385] ? t[166] : t[123];
  assign t[172] = ~(t[164] | t[190]);
  assign t[173] = ~(t[181] | t[177]);
  assign t[174] = ~(t[423]);
  assign t[175] = ~(t[418] | t[419]);
  assign t[176] = ~(t[164] | t[191]);
  assign t[177] = ~(t[164] | t[192]);
  assign t[178] = ~(t[31]);
  assign t[179] = ~(t[424]);
  assign t[17] = ~(t[387] & t[388]);
  assign t[180] = ~(t[421] | t[422]);
  assign t[181] = ~(t[164] | t[193]);
  assign t[182] = ~(t[194] & t[31]);
  assign t[183] = ~(t[164] | t[195]);
  assign t[184] = ~(t[386]);
  assign t[185] = ~(x[7] & t[187]);
  assign t[186] = ~(t[166] & t[185]);
  assign t[187] = ~(t[386] | t[159]);
  assign t[188] = t[164] & t[385];
  assign t[189] = t[385] ? t[196] : t[122];
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = t[385] ? t[197] : t[121];
  assign t[191] = t[385] ? t[123] : t[166];
  assign t[192] = t[385] ? t[122] : t[196];
  assign t[193] = t[385] ? t[185] : t[124];
  assign t[194] = ~(t[172] | t[51]);
  assign t[195] = t[385] ? t[121] : t[197];
  assign t[196] = ~(t[158] & t[388]);
  assign t[197] = ~(t[160] & t[388]);
  assign t[198] = t[1] ? t[199] : t[425];
  assign t[199] = x[6] ? t[201] : t[200];
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = x[7] ? t[203] : t[202];
  assign t[201] = t[204] ^ x[117];
  assign t[202] = t[205] ^ t[206];
  assign t[203] = ~(t[207] ^ t[208]);
  assign t[204] = x[118] ^ x[119];
  assign t[205] = t[30] ? x[119] : x[118];
  assign t[206] = ~(t[209] ^ t[210]);
  assign t[207] = x[7] ? t[212] : t[211];
  assign t[208] = ~(t[213] ^ t[214]);
  assign t[209] = x[7] ? t[216] : t[215];
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = ~(t[217] ^ t[218]);
  assign t[211] = ~(t[219] & t[220]);
  assign t[212] = t[221] ^ t[222];
  assign t[213] = x[7] ? t[224] : t[223];
  assign t[214] = x[7] ? t[226] : t[225];
  assign t[215] = ~(t[227] & t[228]);
  assign t[216] = t[229] ^ t[215];
  assign t[217] = x[7] ? t[231] : t[230];
  assign t[218] = x[7] ? t[233] : t[232];
  assign t[219] = ~(t[391] & t[54]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = ~(t[400] & t[234]);
  assign t[221] = t[91] ? x[121] : x[120];
  assign t[222] = ~(t[235] & t[236]);
  assign t[223] = ~(t[237] & t[238]);
  assign t[224] = t[239] ^ t[232];
  assign t[225] = ~(t[240] & t[241]);
  assign t[226] = t[242] ^ t[223];
  assign t[227] = ~(t[396] & t[67]);
  assign t[228] = ~(t[407] & t[243]);
  assign t[229] = t[30] ? x[123] : x[122];
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = ~(t[244] & t[245]);
  assign t[231] = t[246] ^ t[247];
  assign t[232] = ~(t[248] & t[249]);
  assign t[233] = t[250] ^ t[251];
  assign t[234] = ~(t[392] & t[53]);
  assign t[235] = ~(t[401] & t[89]);
  assign t[236] = ~(t[414] & t[252]);
  assign t[237] = ~(t[405] & t[99]);
  assign t[238] = ~(t[416] & t[253]);
  assign t[239] = t[137] ? x[125] : x[124];
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = ~(t[403] & t[94]);
  assign t[241] = ~(t[415] & t[254]);
  assign t[242] = t[137] ? x[127] : x[126];
  assign t[243] = ~(t[397] & t[66]);
  assign t[244] = ~(t[411] & t[115]);
  assign t[245] = ~(t[420] & t[255]);
  assign t[246] = t[137] ? x[129] : x[128];
  assign t[247] = ~(t[256] & t[257]);
  assign t[248] = ~(t[408] & t[108]);
  assign t[249] = ~(t[417] & t[258]);
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = t[30] ? x[131] : x[130];
  assign t[251] = ~(t[259] & t[260]);
  assign t[252] = ~(t[402] & t[88]);
  assign t[253] = ~(t[406] & t[98]);
  assign t[254] = ~(t[404] & t[93]);
  assign t[255] = ~(t[412] & t[114]);
  assign t[256] = ~(t[421] & t[154]);
  assign t[257] = ~(t[424] & t[261]);
  assign t[258] = ~(t[409] & t[107]);
  assign t[259] = ~(t[418] & t[147]);
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = ~(t[423] & t[262]);
  assign t[261] = ~(t[422] & t[153]);
  assign t[262] = ~(t[419] & t[146]);
  assign t[263] = t[1] ? t[264] : t[426];
  assign t[264] = x[6] ? t[266] : t[265];
  assign t[265] = x[7] ? t[268] : t[267];
  assign t[266] = t[269] ^ x[133];
  assign t[267] = t[270] ^ t[271];
  assign t[268] = ~(t[272] ^ t[273]);
  assign t[269] = x[134] ^ x[135];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[30] ? x[135] : x[134];
  assign t[271] = ~(t[274] ^ t[275]);
  assign t[272] = x[7] ? t[277] : t[276];
  assign t[273] = ~(t[278] ^ t[279]);
  assign t[274] = x[7] ? t[281] : t[280];
  assign t[275] = ~(t[282] ^ t[283]);
  assign t[276] = ~(t[284] & t[285]);
  assign t[277] = t[286] ^ t[287];
  assign t[278] = x[7] ? t[289] : t[288];
  assign t[279] = x[7] ? t[291] : t[290];
  assign t[27] = ~(t[26] ^ t[43]);
  assign t[280] = ~(t[292] & t[293]);
  assign t[281] = t[294] ^ t[280];
  assign t[282] = x[7] ? t[296] : t[295];
  assign t[283] = x[7] ? t[298] : t[297];
  assign t[284] = ~(t[54] & t[86]);
  assign t[285] = ~(t[299] & t[389]);
  assign t[286] = t[91] ? x[137] : x[136];
  assign t[287] = ~(t[300] & t[301]);
  assign t[288] = ~(t[302] & t[303]);
  assign t[289] = t[304] ^ t[290];
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = ~(t[305] & t[306]);
  assign t[291] = t[307] ^ t[297];
  assign t[292] = ~(t[67] & t[103]);
  assign t[293] = ~(t[308] & t[390]);
  assign t[294] = t[30] ? x[139] : x[138];
  assign t[295] = ~(t[309] & t[310]);
  assign t[296] = t[311] ^ t[312];
  assign t[297] = ~(t[313] & t[314]);
  assign t[298] = t[315] ^ t[316];
  assign t[299] = ~(t[317] & t[53]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = ~(t[89] & t[131]);
  assign t[301] = ~(t[318] & t[393]);
  assign t[302] = ~(t[94] & t[135]);
  assign t[303] = ~(t[319] & t[394]);
  assign t[304] = t[137] ? x[141] : x[140];
  assign t[305] = ~(t[99] & t[140]);
  assign t[306] = ~(t[320] & t[395]);
  assign t[307] = t[137] ? x[143] : x[142];
  assign t[308] = ~(t[321] & t[66]);
  assign t[309] = ~(t[115] & t[151]);
  assign t[30] = ~(t[48]);
  assign t[310] = ~(t[322] & t[399]);
  assign t[311] = t[137] ? x[145] : x[144];
  assign t[312] = ~(t[323] & t[324]);
  assign t[313] = ~(t[108] & t[144]);
  assign t[314] = ~(t[325] & t[398]);
  assign t[315] = t[30] ? x[147] : x[146];
  assign t[316] = ~(t[326] & t[327]);
  assign t[317] = ~(t[400] & t[392]);
  assign t[318] = ~(t[328] & t[88]);
  assign t[319] = ~(t[329] & t[93]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = ~(t[330] & t[98]);
  assign t[321] = ~(t[407] & t[397]);
  assign t[322] = ~(t[331] & t[114]);
  assign t[323] = ~(t[154] & t[179]);
  assign t[324] = ~(t[332] & t[413]);
  assign t[325] = ~(t[333] & t[107]);
  assign t[326] = ~(t[147] & t[174]);
  assign t[327] = ~(t[334] & t[410]);
  assign t[328] = ~(t[414] & t[402]);
  assign t[329] = ~(t[415] & t[404]);
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = ~(t[416] & t[406]);
  assign t[331] = ~(t[420] & t[412]);
  assign t[332] = ~(t[335] & t[153]);
  assign t[333] = ~(t[417] & t[409]);
  assign t[334] = ~(t[336] & t[146]);
  assign t[335] = ~(t[424] & t[422]);
  assign t[336] = ~(t[423] & t[419]);
  assign t[337] = t[1] ? t[338] : t[427];
  assign t[338] = x[6] ? t[340] : t[339];
  assign t[339] = x[7] ? t[342] : t[341];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[343] ^ x[149];
  assign t[341] = t[344] ^ t[345];
  assign t[342] = ~(t[346] ^ t[347]);
  assign t[343] = x[150] ^ x[151];
  assign t[344] = t[30] ? x[151] : x[150];
  assign t[345] = ~(t[348] ^ t[349]);
  assign t[346] = x[7] ? t[351] : t[350];
  assign t[347] = ~(t[352] ^ t[353]);
  assign t[348] = x[7] ? t[355] : t[354];
  assign t[349] = ~(t[356] ^ t[357]);
  assign t[34] = ~(t[389] | t[55]);
  assign t[350] = ~(t[284] & t[358]);
  assign t[351] = t[359] ^ t[360];
  assign t[352] = x[7] ? t[362] : t[361];
  assign t[353] = x[7] ? t[364] : t[363];
  assign t[354] = ~(t[292] & t[365]);
  assign t[355] = t[366] ^ t[354];
  assign t[356] = x[7] ? t[368] : t[367];
  assign t[357] = x[7] ? t[370] : t[369];
  assign t[358] = t[33] | t[389];
  assign t[359] = t[91] ? x[153] : x[152];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = ~(t[300] & t[371]);
  assign t[361] = ~(t[302] & t[372]);
  assign t[362] = t[373] ^ t[363];
  assign t[363] = ~(t[305] & t[374]);
  assign t[364] = t[375] ^ t[369];
  assign t[365] = t[41] | t[390];
  assign t[366] = t[30] ? x[155] : x[154];
  assign t[367] = ~(t[309] & t[376]);
  assign t[368] = t[377] ^ t[378];
  assign t[369] = ~(t[313] & t[379]);
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[380] ^ t[381];
  assign t[371] = t[56] | t[393];
  assign t[372] = t[60] | t[394];
  assign t[373] = t[137] ? x[157] : x[156];
  assign t[374] = t[63] | t[395];
  assign t[375] = t[137] ? x[159] : x[158];
  assign t[376] = t[75] | t[399];
  assign t[377] = t[137] ? x[161] : x[160];
  assign t[378] = ~(t[323] & t[382]);
  assign t[379] = t[71] | t[398];
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = t[30] ? x[163] : x[162];
  assign t[381] = ~(t[326] & t[383]);
  assign t[382] = t[117] | t[413];
  assign t[383] = t[110] | t[410];
  assign t[384] = (t[428]);
  assign t[385] = (t[429]);
  assign t[386] = (t[430]);
  assign t[387] = (t[431]);
  assign t[388] = (t[432]);
  assign t[389] = (t[433]);
  assign t[38] = ~(t[39] ^ t[62]);
  assign t[390] = (t[434]);
  assign t[391] = (t[435]);
  assign t[392] = (t[436]);
  assign t[393] = (t[437]);
  assign t[394] = (t[438]);
  assign t[395] = (t[439]);
  assign t[396] = (t[440]);
  assign t[397] = (t[441]);
  assign t[398] = (t[442]);
  assign t[399] = (t[443]);
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (t[444]);
  assign t[401] = (t[445]);
  assign t[402] = (t[446]);
  assign t[403] = (t[447]);
  assign t[404] = (t[448]);
  assign t[405] = (t[449]);
  assign t[406] = (t[450]);
  assign t[407] = (t[451]);
  assign t[408] = (t[452]);
  assign t[409] = (t[453]);
  assign t[40] = ~(t[44] ^ t[65]);
  assign t[410] = (t[454]);
  assign t[411] = (t[455]);
  assign t[412] = (t[456]);
  assign t[413] = (t[457]);
  assign t[414] = (t[458]);
  assign t[415] = (t[459]);
  assign t[416] = (t[460]);
  assign t[417] = (t[461]);
  assign t[418] = (t[462]);
  assign t[419] = (t[463]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (t[464]);
  assign t[421] = (t[465]);
  assign t[422] = (t[466]);
  assign t[423] = (t[467]);
  assign t[424] = (t[468]);
  assign t[425] = (t[469]);
  assign t[426] = (t[470]);
  assign t[427] = (t[471]);
  assign t[428] = t[472] ^ x[5];
  assign t[429] = t[473] ^ x[13];
  assign t[42] = ~(t[390] | t[68]);
  assign t[430] = t[474] ^ x[16];
  assign t[431] = t[475] ^ x[19];
  assign t[432] = t[476] ^ x[22];
  assign t[433] = t[477] ^ x[28];
  assign t[434] = t[478] ^ x[34];
  assign t[435] = t[479] ^ x[35];
  assign t[436] = t[480] ^ x[36];
  assign t[437] = t[481] ^ x[42];
  assign t[438] = t[482] ^ x[50];
  assign t[439] = t[483] ^ x[56];
  assign t[43] = ~(t[69] ^ t[70]);
  assign t[440] = t[484] ^ x[57];
  assign t[441] = t[485] ^ x[58];
  assign t[442] = t[486] ^ x[66];
  assign t[443] = t[487] ^ x[72];
  assign t[444] = t[488] ^ x[73];
  assign t[445] = t[489] ^ x[74];
  assign t[446] = t[490] ^ x[75];
  assign t[447] = t[491] ^ x[76];
  assign t[448] = t[492] ^ x[77];
  assign t[449] = t[493] ^ x[80];
  assign t[44] = ~(t[71] | t[72]);
  assign t[450] = t[494] ^ x[81];
  assign t[451] = t[495] ^ x[84];
  assign t[452] = t[496] ^ x[85];
  assign t[453] = t[497] ^ x[86];
  assign t[454] = t[498] ^ x[92];
  assign t[455] = t[499] ^ x[95];
  assign t[456] = t[500] ^ x[96];
  assign t[457] = t[501] ^ x[102];
  assign t[458] = t[502] ^ x[105];
  assign t[459] = t[503] ^ x[106];
  assign t[45] = ~(t[73] ^ t[74]);
  assign t[460] = t[504] ^ x[107];
  assign t[461] = t[505] ^ x[108];
  assign t[462] = t[506] ^ x[109];
  assign t[463] = t[507] ^ x[110];
  assign t[464] = t[508] ^ x[111];
  assign t[465] = t[509] ^ x[112];
  assign t[466] = t[510] ^ x[113];
  assign t[467] = t[511] ^ x[114];
  assign t[468] = t[512] ^ x[115];
  assign t[469] = t[513] ^ x[116];
  assign t[46] = ~(t[75] | t[76]);
  assign t[470] = t[514] ^ x[132];
  assign t[471] = t[515] ^ x[148];
  assign t[472] = (~t[516] & t[517]);
  assign t[473] = (~t[518] & t[519]);
  assign t[474] = (~t[520] & t[521]);
  assign t[475] = (~t[522] & t[523]);
  assign t[476] = (~t[524] & t[525]);
  assign t[477] = (~t[526] & t[527]);
  assign t[478] = (~t[528] & t[529]);
  assign t[479] = (~t[526] & t[530]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[480] = (~t[526] & t[531]);
  assign t[481] = (~t[532] & t[533]);
  assign t[482] = (~t[534] & t[535]);
  assign t[483] = (~t[536] & t[537]);
  assign t[484] = (~t[528] & t[538]);
  assign t[485] = (~t[528] & t[539]);
  assign t[486] = (~t[540] & t[541]);
  assign t[487] = (~t[542] & t[543]);
  assign t[488] = (~t[526] & t[544]);
  assign t[489] = (~t[532] & t[545]);
  assign t[48] = ~(t[387]);
  assign t[490] = (~t[532] & t[546]);
  assign t[491] = (~t[534] & t[547]);
  assign t[492] = (~t[534] & t[548]);
  assign t[493] = (~t[536] & t[549]);
  assign t[494] = (~t[536] & t[550]);
  assign t[495] = (~t[528] & t[551]);
  assign t[496] = (~t[540] & t[552]);
  assign t[497] = (~t[540] & t[553]);
  assign t[498] = (~t[554] & t[555]);
  assign t[499] = (~t[542] & t[556]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[500] = (~t[542] & t[557]);
  assign t[501] = (~t[558] & t[559]);
  assign t[502] = (~t[532] & t[560]);
  assign t[503] = (~t[534] & t[561]);
  assign t[504] = (~t[536] & t[562]);
  assign t[505] = (~t[540] & t[563]);
  assign t[506] = (~t[554] & t[564]);
  assign t[507] = (~t[554] & t[565]);
  assign t[508] = (~t[542] & t[566]);
  assign t[509] = (~t[558] & t[567]);
  assign t[50] = ~(t[79] | t[81]);
  assign t[510] = (~t[558] & t[568]);
  assign t[511] = (~t[554] & t[569]);
  assign t[512] = (~t[558] & t[570]);
  assign t[513] = (~t[516] & t[571]);
  assign t[514] = (~t[516] & t[572]);
  assign t[515] = (~t[516] & t[573]);
  assign t[516] = t[574] ^ x[4];
  assign t[517] = t[575] ^ x[5];
  assign t[518] = t[576] ^ x[12];
  assign t[519] = t[577] ^ x[13];
  assign t[51] = ~(t[82] & t[83]);
  assign t[520] = t[578] ^ x[15];
  assign t[521] = t[579] ^ x[16];
  assign t[522] = t[580] ^ x[18];
  assign t[523] = t[581] ^ x[19];
  assign t[524] = t[582] ^ x[21];
  assign t[525] = t[583] ^ x[22];
  assign t[526] = t[584] ^ x[27];
  assign t[527] = t[585] ^ x[28];
  assign t[528] = t[586] ^ x[33];
  assign t[529] = t[587] ^ x[34];
  assign t[52] = ~(t[84] & t[85]);
  assign t[530] = t[588] ^ x[35];
  assign t[531] = t[589] ^ x[36];
  assign t[532] = t[590] ^ x[41];
  assign t[533] = t[591] ^ x[42];
  assign t[534] = t[592] ^ x[49];
  assign t[535] = t[593] ^ x[50];
  assign t[536] = t[594] ^ x[55];
  assign t[537] = t[595] ^ x[56];
  assign t[538] = t[596] ^ x[57];
  assign t[539] = t[597] ^ x[58];
  assign t[53] = ~(t[391]);
  assign t[540] = t[598] ^ x[65];
  assign t[541] = t[599] ^ x[66];
  assign t[542] = t[600] ^ x[71];
  assign t[543] = t[601] ^ x[72];
  assign t[544] = t[602] ^ x[73];
  assign t[545] = t[603] ^ x[74];
  assign t[546] = t[604] ^ x[75];
  assign t[547] = t[605] ^ x[76];
  assign t[548] = t[606] ^ x[77];
  assign t[549] = t[607] ^ x[80];
  assign t[54] = ~(t[392]);
  assign t[550] = t[608] ^ x[81];
  assign t[551] = t[609] ^ x[84];
  assign t[552] = t[610] ^ x[85];
  assign t[553] = t[611] ^ x[86];
  assign t[554] = t[612] ^ x[91];
  assign t[555] = t[613] ^ x[92];
  assign t[556] = t[614] ^ x[95];
  assign t[557] = t[615] ^ x[96];
  assign t[558] = t[616] ^ x[101];
  assign t[559] = t[617] ^ x[102];
  assign t[55] = ~(t[86] | t[87]);
  assign t[560] = t[618] ^ x[105];
  assign t[561] = t[619] ^ x[106];
  assign t[562] = t[620] ^ x[107];
  assign t[563] = t[621] ^ x[108];
  assign t[564] = t[622] ^ x[109];
  assign t[565] = t[623] ^ x[110];
  assign t[566] = t[624] ^ x[111];
  assign t[567] = t[625] ^ x[112];
  assign t[568] = t[626] ^ x[113];
  assign t[569] = t[627] ^ x[114];
  assign t[56] = ~(t[88] | t[89]);
  assign t[570] = t[628] ^ x[115];
  assign t[571] = t[629] ^ x[116];
  assign t[572] = t[630] ^ x[132];
  assign t[573] = t[631] ^ x[148];
  assign t[574] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[575] = (x[0]);
  assign t[576] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[577] = (x[11]);
  assign t[578] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[579] = (x[14]);
  assign t[57] = ~(t[393] | t[90]);
  assign t[580] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[581] = (x[17]);
  assign t[582] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[583] = (x[20]);
  assign t[584] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[585] = (x[24]);
  assign t[586] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[587] = (x[30]);
  assign t[588] = (x[25]);
  assign t[589] = (x[26]);
  assign t[58] = t[91] ? x[44] : x[43];
  assign t[590] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[591] = (x[38]);
  assign t[592] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[593] = (x[46]);
  assign t[594] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[595] = (x[52]);
  assign t[596] = (x[31]);
  assign t[597] = (x[32]);
  assign t[598] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[599] = (x[62]);
  assign t[59] = ~(t[92] & t[84]);
  assign t[5] = t[9] ^ x[8];
  assign t[600] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[601] = (x[68]);
  assign t[602] = (x[23]);
  assign t[603] = (x[39]);
  assign t[604] = (x[40]);
  assign t[605] = (x[47]);
  assign t[606] = (x[48]);
  assign t[607] = (x[53]);
  assign t[608] = (x[54]);
  assign t[609] = (x[29]);
  assign t[60] = ~(t[93] | t[94]);
  assign t[610] = (x[63]);
  assign t[611] = (x[64]);
  assign t[612] = (x[87] & ~x[88] & ~x[89] & ~x[90]) | (~x[87] & x[88] & ~x[89] & ~x[90]) | (~x[87] & ~x[88] & x[89] & ~x[90]) | (~x[87] & ~x[88] & ~x[89] & x[90]) | (x[87] & x[88] & x[89] & ~x[90]) | (x[87] & x[88] & ~x[89] & x[90]) | (x[87] & ~x[88] & x[89] & x[90]) | (~x[87] & x[88] & x[89] & x[90]);
  assign t[613] = (x[88]);
  assign t[614] = (x[69]);
  assign t[615] = (x[70]);
  assign t[616] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[617] = (x[98]);
  assign t[618] = (x[37]);
  assign t[619] = (x[45]);
  assign t[61] = ~(t[394] | t[95]);
  assign t[620] = (x[51]);
  assign t[621] = (x[61]);
  assign t[622] = (x[89]);
  assign t[623] = (x[90]);
  assign t[624] = (x[67]);
  assign t[625] = (x[99]);
  assign t[626] = (x[100]);
  assign t[627] = (x[87]);
  assign t[628] = (x[97]);
  assign t[629] = (x[1]);
  assign t[62] = ~(t[96] ^ t[97]);
  assign t[630] = (x[2]);
  assign t[631] = (x[3]);
  assign t[63] = ~(t[98] | t[99]);
  assign t[64] = ~(t[395] | t[100]);
  assign t[65] = ~(t[101] ^ t[102]);
  assign t[66] = ~(t[396]);
  assign t[67] = ~(t[397]);
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = t[30] ? x[60] : x[59];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[107] | t[108]);
  assign t[72] = ~(t[398] | t[109]);
  assign t[73] = ~(t[110] | t[111]);
  assign t[74] = ~(t[112] ^ t[113]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[399] | t[116]);
  assign t[77] = ~(t[117] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[387]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[385] ? t[122] : t[121];
  assign t[81] = t[385] ? t[124] : t[123];
  assign t[82] = ~(t[125] | t[126]);
  assign t[83] = ~(t[79] & t[127]);
  assign t[84] = ~(t[128] & t[129]);
  assign t[85] = t[79] | t[130];
  assign t[86] = ~(t[400]);
  assign t[87] = ~(t[391] | t[392]);
  assign t[88] = ~(t[401]);
  assign t[89] = ~(t[402]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = ~(t[48]);
  assign t[92] = ~(t[133] | t[134]);
  assign t[93] = ~(t[403]);
  assign t[94] = ~(t[404]);
  assign t[95] = ~(t[135] | t[136]);
  assign t[96] = t[137] ? x[79] : x[78];
  assign t[97] = t[138] | t[139];
  assign t[98] = ~(t[405]);
  assign t[99] = ~(t[406]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[198] & ~t[263] & ~t[337]) | (~t[0] & t[198] & ~t[263] & ~t[337]) | (~t[0] & ~t[198] & t[263] & ~t[337]) | (~t[0] & ~t[198] & ~t[263] & t[337]) | (t[0] & t[198] & t[263] & ~t[337]) | (t[0] & t[198] & ~t[263] & t[337]) | (t[0] & ~t[198] & t[263] & t[337]) | (~t[0] & t[198] & t[263] & t[337]);
endmodule

module R2ind181(x, y);
 input [115:0] x;
 output y;

 wire [335:0] t;
  assign t[0] = t[1] ? t[2] : t[103];
  assign t[100] = ~(t[102] | t[98]);
  assign t[101] = ~(t[142]);
  assign t[102] = ~(t[143]);
  assign t[103] = (t[144]);
  assign t[104] = (t[145]);
  assign t[105] = (t[146]);
  assign t[106] = (t[147]);
  assign t[107] = (t[148]);
  assign t[108] = (t[149]);
  assign t[109] = (t[150]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[151]);
  assign t[111] = (t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = t[185] ^ x[5];
  assign t[145] = t[186] ^ x[13];
  assign t[146] = t[187] ^ x[16];
  assign t[147] = t[188] ^ x[19];
  assign t[148] = t[189] ^ x[22];
  assign t[149] = t[190] ^ x[28];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[191] ^ x[36];
  assign t[151] = t[192] ^ x[39];
  assign t[152] = t[193] ^ x[40];
  assign t[153] = t[194] ^ x[46];
  assign t[154] = t[195] ^ x[52];
  assign t[155] = t[196] ^ x[60];
  assign t[156] = t[197] ^ x[63];
  assign t[157] = t[198] ^ x[64];
  assign t[158] = t[199] ^ x[70];
  assign t[159] = t[200] ^ x[78];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[81];
  assign t[161] = t[202] ^ x[82];
  assign t[162] = t[203] ^ x[83];
  assign t[163] = t[204] ^ x[84];
  assign t[164] = t[205] ^ x[85];
  assign t[165] = t[206] ^ x[86];
  assign t[166] = t[207] ^ x[87];
  assign t[167] = t[208] ^ x[88];
  assign t[168] = t[209] ^ x[89];
  assign t[169] = t[210] ^ x[90];
  assign t[16] = ~(t[104] & t[105]);
  assign t[170] = t[211] ^ x[96];
  assign t[171] = t[212] ^ x[97];
  assign t[172] = t[213] ^ x[98];
  assign t[173] = t[214] ^ x[104];
  assign t[174] = t[215] ^ x[105];
  assign t[175] = t[216] ^ x[106];
  assign t[176] = t[217] ^ x[107];
  assign t[177] = t[218] ^ x[108];
  assign t[178] = t[219] ^ x[109];
  assign t[179] = t[220] ^ x[110];
  assign t[17] = ~(t[106] & t[107]);
  assign t[180] = t[221] ^ x[111];
  assign t[181] = t[222] ^ x[112];
  assign t[182] = t[223] ^ x[113];
  assign t[183] = t[224] ^ x[114];
  assign t[184] = t[225] ^ x[115];
  assign t[185] = (~t[226] & t[227]);
  assign t[186] = (~t[228] & t[229]);
  assign t[187] = (~t[230] & t[231]);
  assign t[188] = (~t[232] & t[233]);
  assign t[189] = (~t[234] & t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = (~t[236] & t[237]);
  assign t[191] = (~t[238] & t[239]);
  assign t[192] = (~t[236] & t[240]);
  assign t[193] = (~t[236] & t[241]);
  assign t[194] = (~t[242] & t[243]);
  assign t[195] = (~t[244] & t[245]);
  assign t[196] = (~t[246] & t[247]);
  assign t[197] = (~t[238] & t[248]);
  assign t[198] = (~t[238] & t[249]);
  assign t[199] = (~t[250] & t[251]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[252] & t[253]);
  assign t[201] = (~t[236] & t[254]);
  assign t[202] = (~t[242] & t[255]);
  assign t[203] = (~t[242] & t[256]);
  assign t[204] = (~t[244] & t[257]);
  assign t[205] = (~t[244] & t[258]);
  assign t[206] = (~t[246] & t[259]);
  assign t[207] = (~t[246] & t[260]);
  assign t[208] = (~t[238] & t[261]);
  assign t[209] = (~t[250] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[250] & t[263]);
  assign t[211] = (~t[264] & t[265]);
  assign t[212] = (~t[252] & t[266]);
  assign t[213] = (~t[252] & t[267]);
  assign t[214] = (~t[268] & t[269]);
  assign t[215] = (~t[242] & t[270]);
  assign t[216] = (~t[244] & t[271]);
  assign t[217] = (~t[246] & t[272]);
  assign t[218] = (~t[250] & t[273]);
  assign t[219] = (~t[264] & t[274]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[264] & t[275]);
  assign t[221] = (~t[252] & t[276]);
  assign t[222] = (~t[268] & t[277]);
  assign t[223] = (~t[268] & t[278]);
  assign t[224] = (~t[264] & t[279]);
  assign t[225] = (~t[268] & t[280]);
  assign t[226] = t[281] ^ x[4];
  assign t[227] = t[282] ^ x[5];
  assign t[228] = t[283] ^ x[12];
  assign t[229] = t[284] ^ x[13];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[285] ^ x[15];
  assign t[231] = t[286] ^ x[16];
  assign t[232] = t[287] ^ x[18];
  assign t[233] = t[288] ^ x[19];
  assign t[234] = t[289] ^ x[21];
  assign t[235] = t[290] ^ x[22];
  assign t[236] = t[291] ^ x[27];
  assign t[237] = t[292] ^ x[28];
  assign t[238] = t[293] ^ x[35];
  assign t[239] = t[294] ^ x[36];
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = t[295] ^ x[39];
  assign t[241] = t[296] ^ x[40];
  assign t[242] = t[297] ^ x[45];
  assign t[243] = t[298] ^ x[46];
  assign t[244] = t[299] ^ x[51];
  assign t[245] = t[300] ^ x[52];
  assign t[246] = t[301] ^ x[59];
  assign t[247] = t[302] ^ x[60];
  assign t[248] = t[303] ^ x[63];
  assign t[249] = t[304] ^ x[64];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[305] ^ x[69];
  assign t[251] = t[306] ^ x[70];
  assign t[252] = t[307] ^ x[77];
  assign t[253] = t[308] ^ x[78];
  assign t[254] = t[309] ^ x[81];
  assign t[255] = t[310] ^ x[82];
  assign t[256] = t[311] ^ x[83];
  assign t[257] = t[312] ^ x[84];
  assign t[258] = t[313] ^ x[85];
  assign t[259] = t[314] ^ x[86];
  assign t[25] = ~(t[106]);
  assign t[260] = t[315] ^ x[87];
  assign t[261] = t[316] ^ x[88];
  assign t[262] = t[317] ^ x[89];
  assign t[263] = t[318] ^ x[90];
  assign t[264] = t[319] ^ x[95];
  assign t[265] = t[320] ^ x[96];
  assign t[266] = t[321] ^ x[97];
  assign t[267] = t[322] ^ x[98];
  assign t[268] = t[323] ^ x[103];
  assign t[269] = t[324] ^ x[104];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[325] ^ x[105];
  assign t[271] = t[326] ^ x[106];
  assign t[272] = t[327] ^ x[107];
  assign t[273] = t[328] ^ x[108];
  assign t[274] = t[329] ^ x[109];
  assign t[275] = t[330] ^ x[110];
  assign t[276] = t[331] ^ x[111];
  assign t[277] = t[332] ^ x[112];
  assign t[278] = t[333] ^ x[113];
  assign t[279] = t[334] ^ x[114];
  assign t[27] = t[40] ^ t[26];
  assign t[280] = t[335] ^ x[115];
  assign t[281] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[282] = (x[3]);
  assign t[283] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[284] = (x[11]);
  assign t[285] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[286] = (x[14]);
  assign t[287] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[288] = (x[17]);
  assign t[289] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[290] = (x[20]);
  assign t[291] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[292] = (x[24]);
  assign t[293] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[294] = (x[32]);
  assign t[295] = (x[26]);
  assign t[296] = (x[23]);
  assign t[297] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[298] = (x[42]);
  assign t[299] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[48]);
  assign t[301] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[302] = (x[56]);
  assign t[303] = (x[34]);
  assign t[304] = (x[31]);
  assign t[305] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[306] = (x[66]);
  assign t[307] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[308] = (x[74]);
  assign t[309] = (x[25]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[44]);
  assign t[311] = (x[41]);
  assign t[312] = (x[50]);
  assign t[313] = (x[47]);
  assign t[314] = (x[58]);
  assign t[315] = (x[55]);
  assign t[316] = (x[33]);
  assign t[317] = (x[68]);
  assign t[318] = (x[65]);
  assign t[319] = (x[91] & ~x[92] & ~x[93] & ~x[94]) | (~x[91] & x[92] & ~x[93] & ~x[94]) | (~x[91] & ~x[92] & x[93] & ~x[94]) | (~x[91] & ~x[92] & ~x[93] & x[94]) | (x[91] & x[92] & x[93] & ~x[94]) | (x[91] & x[92] & ~x[93] & x[94]) | (x[91] & ~x[92] & x[93] & x[94]) | (~x[91] & x[92] & x[93] & x[94]);
  assign t[31] = t[47] | t[108];
  assign t[320] = (x[92]);
  assign t[321] = (x[76]);
  assign t[322] = (x[73]);
  assign t[323] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[324] = (x[100]);
  assign t[325] = (x[43]);
  assign t[326] = (x[49]);
  assign t[327] = (x[57]);
  assign t[328] = (x[67]);
  assign t[329] = (x[94]);
  assign t[32] = t[48] ? x[30] : x[29];
  assign t[330] = (x[91]);
  assign t[331] = (x[75]);
  assign t[332] = (x[102]);
  assign t[333] = (x[99]);
  assign t[334] = (x[93]);
  assign t[335] = (x[101]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[36];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[43];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = t[59] | t[109];
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[38] : x[37];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[110]);
  assign t[46] = ~(t[111]);
  assign t[47] = ~(t[68] | t[45]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[69] & t[70]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[71] | t[112];
  assign t[51] = ~(t[72] & t[73]);
  assign t[52] = t[74] | t[113];
  assign t[53] = t[75] ? x[54] : x[53];
  assign t[54] = ~(t[76] & t[77]);
  assign t[55] = t[78] | t[114];
  assign t[56] = t[75] ? x[62] : x[61];
  assign t[57] = ~(t[115]);
  assign t[58] = ~(t[116]);
  assign t[59] = ~(t[79] | t[57]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[80] & t[81]);
  assign t[61] = t[82] | t[117];
  assign t[62] = t[75] ? x[72] : x[71];
  assign t[63] = ~(t[83] & t[84]);
  assign t[64] = ~(t[85] & t[86]);
  assign t[65] = t[87] | t[118];
  assign t[66] = t[18] ? x[80] : x[79];
  assign t[67] = ~(t[88] & t[89]);
  assign t[68] = ~(t[119]);
  assign t[69] = ~(t[120]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[121]);
  assign t[71] = ~(t[90] | t[69]);
  assign t[72] = ~(t[122]);
  assign t[73] = ~(t[123]);
  assign t[74] = ~(t[91] | t[72]);
  assign t[75] = ~(t[25]);
  assign t[76] = ~(t[124]);
  assign t[77] = ~(t[125]);
  assign t[78] = ~(t[92] | t[76]);
  assign t[79] = ~(t[126]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[127]);
  assign t[81] = ~(t[128]);
  assign t[82] = ~(t[93] | t[80]);
  assign t[83] = ~(t[94] & t[95]);
  assign t[84] = t[96] | t[129];
  assign t[85] = ~(t[130]);
  assign t[86] = ~(t[131]);
  assign t[87] = ~(t[97] | t[85]);
  assign t[88] = ~(t[98] & t[99]);
  assign t[89] = t[100] | t[132];
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[133]);
  assign t[91] = ~(t[134]);
  assign t[92] = ~(t[135]);
  assign t[93] = ~(t[136]);
  assign t[94] = ~(t[137]);
  assign t[95] = ~(t[138]);
  assign t[96] = ~(t[101] | t[94]);
  assign t[97] = ~(t[139]);
  assign t[98] = ~(t[140]);
  assign t[99] = ~(t[141]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [115:0] x;
 output y;

 wire [344:0] t;
  assign t[0] = t[1] ? t[2] : t[112];
  assign t[100] = ~(t[146]);
  assign t[101] = ~(t[147]);
  assign t[102] = ~(t[108] & t[109]);
  assign t[103] = ~(t[140] & t[139]);
  assign t[104] = ~(t[148]);
  assign t[105] = ~(t[149]);
  assign t[106] = ~(t[150]);
  assign t[107] = ~(t[110] & t[111]);
  assign t[108] = ~(t[147] & t[146]);
  assign t[109] = ~(t[151]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[150] & t[149]);
  assign t[111] = ~(t[152]);
  assign t[112] = (t[153]);
  assign t[113] = (t[154]);
  assign t[114] = (t[155]);
  assign t[115] = (t[156]);
  assign t[116] = (t[157]);
  assign t[117] = (t[158]);
  assign t[118] = (t[159]);
  assign t[119] = (t[160]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[161]);
  assign t[121] = (t[162]);
  assign t[122] = (t[163]);
  assign t[123] = (t[164]);
  assign t[124] = (t[165]);
  assign t[125] = (t[166]);
  assign t[126] = (t[167]);
  assign t[127] = (t[168]);
  assign t[128] = (t[169]);
  assign t[129] = (t[170]);
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = (t[171]);
  assign t[131] = (t[172]);
  assign t[132] = (t[173]);
  assign t[133] = (t[174]);
  assign t[134] = (t[175]);
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = t[194] ^ x[5];
  assign t[154] = t[195] ^ x[13];
  assign t[155] = t[196] ^ x[16];
  assign t[156] = t[197] ^ x[19];
  assign t[157] = t[198] ^ x[22];
  assign t[158] = t[199] ^ x[28];
  assign t[159] = t[200] ^ x[36];
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = t[201] ^ x[39];
  assign t[161] = t[202] ^ x[40];
  assign t[162] = t[203] ^ x[46];
  assign t[163] = t[204] ^ x[52];
  assign t[164] = t[205] ^ x[60];
  assign t[165] = t[206] ^ x[63];
  assign t[166] = t[207] ^ x[64];
  assign t[167] = t[208] ^ x[70];
  assign t[168] = t[209] ^ x[78];
  assign t[169] = t[210] ^ x[81];
  assign t[16] = ~(t[113] & t[114]);
  assign t[170] = t[211] ^ x[82];
  assign t[171] = t[212] ^ x[83];
  assign t[172] = t[213] ^ x[84];
  assign t[173] = t[214] ^ x[85];
  assign t[174] = t[215] ^ x[86];
  assign t[175] = t[216] ^ x[87];
  assign t[176] = t[217] ^ x[88];
  assign t[177] = t[218] ^ x[89];
  assign t[178] = t[219] ^ x[90];
  assign t[179] = t[220] ^ x[96];
  assign t[17] = ~(t[115] & t[116]);
  assign t[180] = t[221] ^ x[97];
  assign t[181] = t[222] ^ x[98];
  assign t[182] = t[223] ^ x[104];
  assign t[183] = t[224] ^ x[105];
  assign t[184] = t[225] ^ x[106];
  assign t[185] = t[226] ^ x[107];
  assign t[186] = t[227] ^ x[108];
  assign t[187] = t[228] ^ x[109];
  assign t[188] = t[229] ^ x[110];
  assign t[189] = t[230] ^ x[111];
  assign t[18] = ~(t[25]);
  assign t[190] = t[231] ^ x[112];
  assign t[191] = t[232] ^ x[113];
  assign t[192] = t[233] ^ x[114];
  assign t[193] = t[234] ^ x[115];
  assign t[194] = (~t[235] & t[236]);
  assign t[195] = (~t[237] & t[238]);
  assign t[196] = (~t[239] & t[240]);
  assign t[197] = (~t[241] & t[242]);
  assign t[198] = (~t[243] & t[244]);
  assign t[199] = (~t[245] & t[246]);
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (~t[247] & t[248]);
  assign t[201] = (~t[245] & t[249]);
  assign t[202] = (~t[245] & t[250]);
  assign t[203] = (~t[251] & t[252]);
  assign t[204] = (~t[253] & t[254]);
  assign t[205] = (~t[255] & t[256]);
  assign t[206] = (~t[247] & t[257]);
  assign t[207] = (~t[247] & t[258]);
  assign t[208] = (~t[259] & t[260]);
  assign t[209] = (~t[261] & t[262]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[245] & t[263]);
  assign t[211] = (~t[251] & t[264]);
  assign t[212] = (~t[251] & t[265]);
  assign t[213] = (~t[253] & t[266]);
  assign t[214] = (~t[253] & t[267]);
  assign t[215] = (~t[255] & t[268]);
  assign t[216] = (~t[255] & t[269]);
  assign t[217] = (~t[247] & t[270]);
  assign t[218] = (~t[259] & t[271]);
  assign t[219] = (~t[259] & t[272]);
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = (~t[273] & t[274]);
  assign t[221] = (~t[261] & t[275]);
  assign t[222] = (~t[261] & t[276]);
  assign t[223] = (~t[277] & t[278]);
  assign t[224] = (~t[251] & t[279]);
  assign t[225] = (~t[253] & t[280]);
  assign t[226] = (~t[255] & t[281]);
  assign t[227] = (~t[259] & t[282]);
  assign t[228] = (~t[273] & t[283]);
  assign t[229] = (~t[273] & t[284]);
  assign t[22] = t[32] ^ t[33];
  assign t[230] = (~t[261] & t[285]);
  assign t[231] = (~t[277] & t[286]);
  assign t[232] = (~t[277] & t[287]);
  assign t[233] = (~t[273] & t[288]);
  assign t[234] = (~t[277] & t[289]);
  assign t[235] = t[290] ^ x[4];
  assign t[236] = t[291] ^ x[5];
  assign t[237] = t[292] ^ x[12];
  assign t[238] = t[293] ^ x[13];
  assign t[239] = t[294] ^ x[15];
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = t[295] ^ x[16];
  assign t[241] = t[296] ^ x[18];
  assign t[242] = t[297] ^ x[19];
  assign t[243] = t[298] ^ x[21];
  assign t[244] = t[299] ^ x[22];
  assign t[245] = t[300] ^ x[27];
  assign t[246] = t[301] ^ x[28];
  assign t[247] = t[302] ^ x[35];
  assign t[248] = t[303] ^ x[36];
  assign t[249] = t[304] ^ x[39];
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = t[305] ^ x[40];
  assign t[251] = t[306] ^ x[45];
  assign t[252] = t[307] ^ x[46];
  assign t[253] = t[308] ^ x[51];
  assign t[254] = t[309] ^ x[52];
  assign t[255] = t[310] ^ x[59];
  assign t[256] = t[311] ^ x[60];
  assign t[257] = t[312] ^ x[63];
  assign t[258] = t[313] ^ x[64];
  assign t[259] = t[314] ^ x[69];
  assign t[25] = ~(t[115]);
  assign t[260] = t[315] ^ x[70];
  assign t[261] = t[316] ^ x[77];
  assign t[262] = t[317] ^ x[78];
  assign t[263] = t[318] ^ x[81];
  assign t[264] = t[319] ^ x[82];
  assign t[265] = t[320] ^ x[83];
  assign t[266] = t[321] ^ x[84];
  assign t[267] = t[322] ^ x[85];
  assign t[268] = t[323] ^ x[86];
  assign t[269] = t[324] ^ x[87];
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = t[325] ^ x[88];
  assign t[271] = t[326] ^ x[89];
  assign t[272] = t[327] ^ x[90];
  assign t[273] = t[328] ^ x[95];
  assign t[274] = t[329] ^ x[96];
  assign t[275] = t[330] ^ x[97];
  assign t[276] = t[331] ^ x[98];
  assign t[277] = t[332] ^ x[103];
  assign t[278] = t[333] ^ x[104];
  assign t[279] = t[334] ^ x[105];
  assign t[27] = t[40] ^ t[26];
  assign t[280] = t[335] ^ x[106];
  assign t[281] = t[336] ^ x[107];
  assign t[282] = t[337] ^ x[108];
  assign t[283] = t[338] ^ x[109];
  assign t[284] = t[339] ^ x[110];
  assign t[285] = t[340] ^ x[111];
  assign t[286] = t[341] ^ x[112];
  assign t[287] = t[342] ^ x[113];
  assign t[288] = t[343] ^ x[114];
  assign t[289] = t[344] ^ x[115];
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[290] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[291] = (x[2]);
  assign t[292] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[293] = (x[11]);
  assign t[294] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[295] = (x[14]);
  assign t[296] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[297] = (x[17]);
  assign t[298] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[299] = (x[20]);
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[301] = (x[24]);
  assign t[302] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[303] = (x[32]);
  assign t[304] = (x[26]);
  assign t[305] = (x[23]);
  assign t[306] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[307] = (x[42]);
  assign t[308] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[309] = (x[48]);
  assign t[30] = ~(t[45] & t[46]);
  assign t[310] = (x[55] & ~x[56] & ~x[57] & ~x[58]) | (~x[55] & x[56] & ~x[57] & ~x[58]) | (~x[55] & ~x[56] & x[57] & ~x[58]) | (~x[55] & ~x[56] & ~x[57] & x[58]) | (x[55] & x[56] & x[57] & ~x[58]) | (x[55] & x[56] & ~x[57] & x[58]) | (x[55] & ~x[56] & x[57] & x[58]) | (~x[55] & x[56] & x[57] & x[58]);
  assign t[311] = (x[56]);
  assign t[312] = (x[34]);
  assign t[313] = (x[31]);
  assign t[314] = (x[65] & ~x[66] & ~x[67] & ~x[68]) | (~x[65] & x[66] & ~x[67] & ~x[68]) | (~x[65] & ~x[66] & x[67] & ~x[68]) | (~x[65] & ~x[66] & ~x[67] & x[68]) | (x[65] & x[66] & x[67] & ~x[68]) | (x[65] & x[66] & ~x[67] & x[68]) | (x[65] & ~x[66] & x[67] & x[68]) | (~x[65] & x[66] & x[67] & x[68]);
  assign t[315] = (x[66]);
  assign t[316] = (x[73] & ~x[74] & ~x[75] & ~x[76]) | (~x[73] & x[74] & ~x[75] & ~x[76]) | (~x[73] & ~x[74] & x[75] & ~x[76]) | (~x[73] & ~x[74] & ~x[75] & x[76]) | (x[73] & x[74] & x[75] & ~x[76]) | (x[73] & x[74] & ~x[75] & x[76]) | (x[73] & ~x[74] & x[75] & x[76]) | (~x[73] & x[74] & x[75] & x[76]);
  assign t[317] = (x[74]);
  assign t[318] = (x[25]);
  assign t[319] = (x[44]);
  assign t[31] = ~(t[47] & t[117]);
  assign t[320] = (x[41]);
  assign t[321] = (x[50]);
  assign t[322] = (x[47]);
  assign t[323] = (x[58]);
  assign t[324] = (x[55]);
  assign t[325] = (x[33]);
  assign t[326] = (x[68]);
  assign t[327] = (x[65]);
  assign t[328] = (x[91] & ~x[92] & ~x[93] & ~x[94]) | (~x[91] & x[92] & ~x[93] & ~x[94]) | (~x[91] & ~x[92] & x[93] & ~x[94]) | (~x[91] & ~x[92] & ~x[93] & x[94]) | (x[91] & x[92] & x[93] & ~x[94]) | (x[91] & x[92] & ~x[93] & x[94]) | (x[91] & ~x[92] & x[93] & x[94]) | (~x[91] & x[92] & x[93] & x[94]);
  assign t[329] = (x[92]);
  assign t[32] = t[48] ? x[30] : x[29];
  assign t[330] = (x[76]);
  assign t[331] = (x[73]);
  assign t[332] = (x[99] & ~x[100] & ~x[101] & ~x[102]) | (~x[99] & x[100] & ~x[101] & ~x[102]) | (~x[99] & ~x[100] & x[101] & ~x[102]) | (~x[99] & ~x[100] & ~x[101] & x[102]) | (x[99] & x[100] & x[101] & ~x[102]) | (x[99] & x[100] & ~x[101] & x[102]) | (x[99] & ~x[100] & x[101] & x[102]) | (~x[99] & x[100] & x[101] & x[102]);
  assign t[333] = (x[100]);
  assign t[334] = (x[43]);
  assign t[335] = (x[49]);
  assign t[336] = (x[57]);
  assign t[337] = (x[67]);
  assign t[338] = (x[94]);
  assign t[339] = (x[91]);
  assign t[33] = ~(t[49] & t[50]);
  assign t[340] = (x[75]);
  assign t[341] = (x[102]);
  assign t[342] = (x[99]);
  assign t[343] = (x[93]);
  assign t[344] = (x[101]);
  assign t[34] = ~(t[51] & t[52]);
  assign t[35] = t[53] ^ t[36];
  assign t[36] = ~(t[54] & t[55]);
  assign t[37] = t[56] ^ t[43];
  assign t[38] = ~(t[57] & t[58]);
  assign t[39] = ~(t[59] & t[118]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[38] : x[37];
  assign t[41] = ~(t[60] & t[61]);
  assign t[42] = t[62] ^ t[63];
  assign t[43] = ~(t[64] & t[65]);
  assign t[44] = t[66] ^ t[67];
  assign t[45] = ~(t[119]);
  assign t[46] = ~(t[120]);
  assign t[47] = ~(t[68] & t[69]);
  assign t[48] = ~(t[25]);
  assign t[49] = ~(t[70] & t[71]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[72] & t[121]);
  assign t[51] = ~(t[73] & t[74]);
  assign t[52] = ~(t[75] & t[122]);
  assign t[53] = t[76] ? x[54] : x[53];
  assign t[54] = ~(t[77] & t[78]);
  assign t[55] = ~(t[79] & t[123]);
  assign t[56] = t[76] ? x[62] : x[61];
  assign t[57] = ~(t[124]);
  assign t[58] = ~(t[125]);
  assign t[59] = ~(t[80] & t[81]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[82] & t[83]);
  assign t[61] = ~(t[84] & t[126]);
  assign t[62] = t[76] ? x[72] : x[71];
  assign t[63] = ~(t[85] & t[86]);
  assign t[64] = ~(t[87] & t[88]);
  assign t[65] = ~(t[89] & t[127]);
  assign t[66] = t[18] ? x[80] : x[79];
  assign t[67] = ~(t[90] & t[91]);
  assign t[68] = ~(t[120] & t[119]);
  assign t[69] = ~(t[128]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[129]);
  assign t[71] = ~(t[130]);
  assign t[72] = ~(t[92] & t[93]);
  assign t[73] = ~(t[131]);
  assign t[74] = ~(t[132]);
  assign t[75] = ~(t[94] & t[95]);
  assign t[76] = ~(t[25]);
  assign t[77] = ~(t[133]);
  assign t[78] = ~(t[134]);
  assign t[79] = ~(t[96] & t[97]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[125] & t[124]);
  assign t[81] = ~(t[135]);
  assign t[82] = ~(t[136]);
  assign t[83] = ~(t[137]);
  assign t[84] = ~(t[98] & t[99]);
  assign t[85] = ~(t[100] & t[101]);
  assign t[86] = ~(t[102] & t[138]);
  assign t[87] = ~(t[139]);
  assign t[88] = ~(t[140]);
  assign t[89] = ~(t[103] & t[104]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[105] & t[106]);
  assign t[91] = ~(t[107] & t[141]);
  assign t[92] = ~(t[130] & t[129]);
  assign t[93] = ~(t[142]);
  assign t[94] = ~(t[132] & t[131]);
  assign t[95] = ~(t[143]);
  assign t[96] = ~(t[134] & t[133]);
  assign t[97] = ~(t[144]);
  assign t[98] = ~(t[137] & t[136]);
  assign t[99] = ~(t[145]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [106:0] x;
 output y;

 wire [281:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[5];
  assign t[127] = t[159] ^ x[13];
  assign t[128] = t[160] ^ x[16];
  assign t[129] = t[161] ^ x[19];
  assign t[12] = t[18] ? x[10] : x[9];
  assign t[130] = t[162] ^ x[22];
  assign t[131] = t[163] ^ x[28];
  assign t[132] = t[164] ^ x[29];
  assign t[133] = t[165] ^ x[37];
  assign t[134] = t[166] ^ x[38];
  assign t[135] = t[167] ^ x[41];
  assign t[136] = t[168] ^ x[47];
  assign t[137] = t[169] ^ x[48];
  assign t[138] = t[170] ^ x[54];
  assign t[139] = t[171] ^ x[55];
  assign t[13] = ~(t[19] ^ t[20]);
  assign t[140] = t[172] ^ x[63];
  assign t[141] = t[173] ^ x[64];
  assign t[142] = t[174] ^ x[67];
  assign t[143] = t[175] ^ x[73];
  assign t[144] = t[176] ^ x[74];
  assign t[145] = t[177] ^ x[82];
  assign t[146] = t[178] ^ x[83];
  assign t[147] = t[179] ^ x[86];
  assign t[148] = t[180] ^ x[87];
  assign t[149] = t[181] ^ x[88];
  assign t[14] = x[7] ? t[22] : t[21];
  assign t[150] = t[182] ^ x[89];
  assign t[151] = t[183] ^ x[95];
  assign t[152] = t[184] ^ x[96];
  assign t[153] = t[185] ^ x[97];
  assign t[154] = t[186] ^ x[103];
  assign t[155] = t[187] ^ x[104];
  assign t[156] = t[188] ^ x[105];
  assign t[157] = t[189] ^ x[106];
  assign t[158] = (~t[190] & t[191]);
  assign t[159] = (~t[192] & t[193]);
  assign t[15] = ~(t[23] ^ t[24]);
  assign t[160] = (~t[194] & t[195]);
  assign t[161] = (~t[196] & t[197]);
  assign t[162] = (~t[198] & t[199]);
  assign t[163] = (~t[200] & t[201]);
  assign t[164] = (~t[200] & t[202]);
  assign t[165] = (~t[203] & t[204]);
  assign t[166] = (~t[203] & t[205]);
  assign t[167] = (~t[200] & t[206]);
  assign t[168] = (~t[207] & t[208]);
  assign t[169] = (~t[207] & t[209]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (~t[210] & t[211]);
  assign t[171] = (~t[210] & t[212]);
  assign t[172] = (~t[213] & t[214]);
  assign t[173] = (~t[213] & t[215]);
  assign t[174] = (~t[203] & t[216]);
  assign t[175] = (~t[217] & t[218]);
  assign t[176] = (~t[217] & t[219]);
  assign t[177] = (~t[220] & t[221]);
  assign t[178] = (~t[220] & t[222]);
  assign t[179] = (~t[207] & t[223]);
  assign t[17] = ~(t[97] & t[98]);
  assign t[180] = (~t[210] & t[224]);
  assign t[181] = (~t[213] & t[225]);
  assign t[182] = (~t[217] & t[226]);
  assign t[183] = (~t[227] & t[228]);
  assign t[184] = (~t[227] & t[229]);
  assign t[185] = (~t[220] & t[230]);
  assign t[186] = (~t[231] & t[232]);
  assign t[187] = (~t[231] & t[233]);
  assign t[188] = (~t[227] & t[234]);
  assign t[189] = (~t[231] & t[235]);
  assign t[18] = ~(t[25]);
  assign t[190] = t[236] ^ x[4];
  assign t[191] = t[237] ^ x[5];
  assign t[192] = t[238] ^ x[12];
  assign t[193] = t[239] ^ x[13];
  assign t[194] = t[240] ^ x[15];
  assign t[195] = t[241] ^ x[16];
  assign t[196] = t[242] ^ x[18];
  assign t[197] = t[243] ^ x[19];
  assign t[198] = t[244] ^ x[21];
  assign t[199] = t[245] ^ x[22];
  assign t[19] = x[7] ? t[27] : t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[246] ^ x[27];
  assign t[201] = t[247] ^ x[28];
  assign t[202] = t[248] ^ x[29];
  assign t[203] = t[249] ^ x[36];
  assign t[204] = t[250] ^ x[37];
  assign t[205] = t[251] ^ x[38];
  assign t[206] = t[252] ^ x[41];
  assign t[207] = t[253] ^ x[46];
  assign t[208] = t[254] ^ x[47];
  assign t[209] = t[255] ^ x[48];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[256] ^ x[53];
  assign t[211] = t[257] ^ x[54];
  assign t[212] = t[258] ^ x[55];
  assign t[213] = t[259] ^ x[62];
  assign t[214] = t[260] ^ x[63];
  assign t[215] = t[261] ^ x[64];
  assign t[216] = t[262] ^ x[67];
  assign t[217] = t[263] ^ x[72];
  assign t[218] = t[264] ^ x[73];
  assign t[219] = t[265] ^ x[74];
  assign t[21] = ~(t[30] & t[31]);
  assign t[220] = t[266] ^ x[81];
  assign t[221] = t[267] ^ x[82];
  assign t[222] = t[268] ^ x[83];
  assign t[223] = t[269] ^ x[86];
  assign t[224] = t[270] ^ x[87];
  assign t[225] = t[271] ^ x[88];
  assign t[226] = t[272] ^ x[89];
  assign t[227] = t[273] ^ x[94];
  assign t[228] = t[274] ^ x[95];
  assign t[229] = t[275] ^ x[96];
  assign t[22] = t[32] ^ t[33];
  assign t[230] = t[276] ^ x[97];
  assign t[231] = t[277] ^ x[102];
  assign t[232] = t[278] ^ x[103];
  assign t[233] = t[279] ^ x[104];
  assign t[234] = t[280] ^ x[105];
  assign t[235] = t[281] ^ x[106];
  assign t[236] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[237] = (x[1]);
  assign t[238] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[239] = (x[11]);
  assign t[23] = x[7] ? t[35] : t[34];
  assign t[240] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[241] = (x[14]);
  assign t[242] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[243] = (x[17]);
  assign t[244] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[245] = (x[20]);
  assign t[246] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[247] = (x[25]);
  assign t[248] = (x[23]);
  assign t[249] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[24] = x[7] ? t[37] : t[36];
  assign t[250] = (x[34]);
  assign t[251] = (x[32]);
  assign t[252] = (x[26]);
  assign t[253] = (x[42] & ~x[43] & ~x[44] & ~x[45]) | (~x[42] & x[43] & ~x[44] & ~x[45]) | (~x[42] & ~x[43] & x[44] & ~x[45]) | (~x[42] & ~x[43] & ~x[44] & x[45]) | (x[42] & x[43] & x[44] & ~x[45]) | (x[42] & x[43] & ~x[44] & x[45]) | (x[42] & ~x[43] & x[44] & x[45]) | (~x[42] & x[43] & x[44] & x[45]);
  assign t[254] = (x[44]);
  assign t[255] = (x[42]);
  assign t[256] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[257] = (x[51]);
  assign t[258] = (x[49]);
  assign t[259] = (x[58] & ~x[59] & ~x[60] & ~x[61]) | (~x[58] & x[59] & ~x[60] & ~x[61]) | (~x[58] & ~x[59] & x[60] & ~x[61]) | (~x[58] & ~x[59] & ~x[60] & x[61]) | (x[58] & x[59] & x[60] & ~x[61]) | (x[58] & x[59] & ~x[60] & x[61]) | (x[58] & ~x[59] & x[60] & x[61]) | (~x[58] & x[59] & x[60] & x[61]);
  assign t[25] = ~(t[97]);
  assign t[260] = (x[60]);
  assign t[261] = (x[58]);
  assign t[262] = (x[35]);
  assign t[263] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[264] = (x[70]);
  assign t[265] = (x[68]);
  assign t[266] = (x[77] & ~x[78] & ~x[79] & ~x[80]) | (~x[77] & x[78] & ~x[79] & ~x[80]) | (~x[77] & ~x[78] & x[79] & ~x[80]) | (~x[77] & ~x[78] & ~x[79] & x[80]) | (x[77] & x[78] & x[79] & ~x[80]) | (x[77] & x[78] & ~x[79] & x[80]) | (x[77] & ~x[78] & x[79] & x[80]) | (~x[77] & x[78] & x[79] & x[80]);
  assign t[267] = (x[79]);
  assign t[268] = (x[77]);
  assign t[269] = (x[45]);
  assign t[26] = ~(t[38] & t[39]);
  assign t[270] = (x[52]);
  assign t[271] = (x[61]);
  assign t[272] = (x[71]);
  assign t[273] = (x[90] & ~x[91] & ~x[92] & ~x[93]) | (~x[90] & x[91] & ~x[92] & ~x[93]) | (~x[90] & ~x[91] & x[92] & ~x[93]) | (~x[90] & ~x[91] & ~x[92] & x[93]) | (x[90] & x[91] & x[92] & ~x[93]) | (x[90] & x[91] & ~x[92] & x[93]) | (x[90] & ~x[91] & x[92] & x[93]) | (~x[90] & x[91] & x[92] & x[93]);
  assign t[274] = (x[92]);
  assign t[275] = (x[90]);
  assign t[276] = (x[80]);
  assign t[277] = (x[98] & ~x[99] & ~x[100] & ~x[101]) | (~x[98] & x[99] & ~x[100] & ~x[101]) | (~x[98] & ~x[99] & x[100] & ~x[101]) | (~x[98] & ~x[99] & ~x[100] & x[101]) | (x[98] & x[99] & x[100] & ~x[101]) | (x[98] & x[99] & ~x[100] & x[101]) | (x[98] & ~x[99] & x[100] & x[101]) | (~x[98] & x[99] & x[100] & x[101]);
  assign t[278] = (x[100]);
  assign t[279] = (x[98]);
  assign t[27] = t[40] ^ t[26];
  assign t[280] = (x[93]);
  assign t[281] = (x[101]);
  assign t[28] = x[7] ? t[42] : t[41];
  assign t[29] = x[7] ? t[44] : t[43];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[99] & t[45]);
  assign t[31] = ~(t[100] & t[46]);
  assign t[32] = t[47] ? x[31] : x[30];
  assign t[33] = ~(t[48] & t[49]);
  assign t[34] = ~(t[50] & t[51]);
  assign t[35] = t[52] ^ t[43];
  assign t[36] = ~(t[53] & t[54]);
  assign t[37] = t[55] ^ t[34];
  assign t[38] = ~(t[101] & t[56]);
  assign t[39] = ~(t[102] & t[57]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[18] ? x[40] : x[39];
  assign t[41] = ~(t[58] & t[59]);
  assign t[42] = t[60] ^ t[61];
  assign t[43] = ~(t[62] & t[63]);
  assign t[44] = t[64] ^ t[65];
  assign t[45] = ~(t[103]);
  assign t[46] = ~(t[103] & t[66]);
  assign t[47] = ~(t[25]);
  assign t[48] = ~(t[104] & t[67]);
  assign t[49] = ~(t[105] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[106] & t[69]);
  assign t[51] = ~(t[107] & t[70]);
  assign t[52] = t[71] ? x[57] : x[56];
  assign t[53] = ~(t[108] & t[72]);
  assign t[54] = ~(t[109] & t[73]);
  assign t[55] = t[71] ? x[66] : x[65];
  assign t[56] = ~(t[110]);
  assign t[57] = ~(t[110] & t[74]);
  assign t[58] = ~(t[111] & t[75]);
  assign t[59] = ~(t[112] & t[76]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[71] ? x[76] : x[75];
  assign t[61] = ~(t[77] & t[78]);
  assign t[62] = ~(t[113] & t[79]);
  assign t[63] = ~(t[114] & t[80]);
  assign t[64] = t[18] ? x[85] : x[84];
  assign t[65] = ~(t[81] & t[82]);
  assign t[66] = ~(t[99]);
  assign t[67] = ~(t[115]);
  assign t[68] = ~(t[115] & t[83]);
  assign t[69] = ~(t[116]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[116] & t[84]);
  assign t[71] = ~(t[25]);
  assign t[72] = ~(t[117]);
  assign t[73] = ~(t[117] & t[85]);
  assign t[74] = ~(t[101]);
  assign t[75] = ~(t[118]);
  assign t[76] = ~(t[118] & t[86]);
  assign t[77] = ~(t[119] & t[87]);
  assign t[78] = ~(t[120] & t[88]);
  assign t[79] = ~(t[121]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[121] & t[89]);
  assign t[81] = ~(t[122] & t[90]);
  assign t[82] = ~(t[123] & t[91]);
  assign t[83] = ~(t[104]);
  assign t[84] = ~(t[106]);
  assign t[85] = ~(t[108]);
  assign t[86] = ~(t[111]);
  assign t[87] = ~(t[124]);
  assign t[88] = ~(t[124] & t[92]);
  assign t[89] = ~(t[113]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[125]);
  assign t[91] = ~(t[125] & t[93]);
  assign t[92] = ~(t[119]);
  assign t[93] = ~(t[122]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [115:0] x;
 output y;

 wire [430:0] t;
  assign t[0] = t[1] ? t[2] : t[198];
  assign t[100] = ~(t[140] | t[141]);
  assign t[101] = t[137] ? x[83] : x[82];
  assign t[102] = ~(t[142] & t[106]);
  assign t[103] = ~(t[221]);
  assign t[104] = ~(t[210] | t[211]);
  assign t[105] = ~(t[125] | t[50]);
  assign t[106] = ~(t[143] | t[139]);
  assign t[107] = ~(t[222]);
  assign t[108] = ~(t[223]);
  assign t[109] = ~(t[144] | t[145]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[110] = ~(t[146] | t[147]);
  assign t[111] = ~(t[224] | t[148]);
  assign t[112] = t[30] ? x[94] : x[93];
  assign t[113] = ~(t[149] & t[150]);
  assign t[114] = ~(t[225]);
  assign t[115] = ~(t[226]);
  assign t[116] = ~(t[151] | t[152]);
  assign t[117] = ~(t[153] | t[154]);
  assign t[118] = ~(t[227] | t[155]);
  assign t[119] = t[137] ? x[104] : x[103];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[156] & t[157]);
  assign t[121] = ~(t[158] & t[159]);
  assign t[122] = ~(t[160] & t[159]);
  assign t[123] = ~(x[7] & t[161]);
  assign t[124] = ~(t[162] & t[159]);
  assign t[125] = ~(t[79] | t[163]);
  assign t[126] = ~(t[164] | t[165]);
  assign t[127] = ~(t[123] & t[166]);
  assign t[128] = t[202] & t[167];
  assign t[129] = t[158] | t[160];
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = t[199] ? t[123] : t[124];
  assign t[131] = ~(t[228]);
  assign t[132] = ~(t[215] | t[216]);
  assign t[133] = ~(t[168] & t[169]);
  assign t[134] = t[139] | t[170];
  assign t[135] = ~(t[229]);
  assign t[136] = ~(t[217] | t[218]);
  assign t[137] = ~(t[48]);
  assign t[138] = ~(t[31] & t[169]);
  assign t[139] = ~(t[164] | t[171]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[140] = ~(t[230]);
  assign t[141] = ~(t[219] | t[220]);
  assign t[142] = ~(t[172]);
  assign t[143] = ~(t[173]);
  assign t[144] = ~(t[231]);
  assign t[145] = ~(t[222] | t[223]);
  assign t[146] = ~(t[232]);
  assign t[147] = ~(t[233]);
  assign t[148] = ~(t[174] | t[175]);
  assign t[149] = ~(t[176] | t[177]);
  assign t[14] = x[7] ? t[23] : t[22];
  assign t[150] = ~(t[128] | t[178]);
  assign t[151] = ~(t[234]);
  assign t[152] = ~(t[225] | t[226]);
  assign t[153] = ~(t[235]);
  assign t[154] = ~(t[236]);
  assign t[155] = ~(t[179] | t[180]);
  assign t[156] = ~(t[181] | t[182]);
  assign t[157] = ~(t[183]);
  assign t[158] = ~(x[7] | t[200]);
  assign t[159] = ~(t[202]);
  assign t[15] = ~(t[24] ^ t[25]);
  assign t[160] = x[7] & t[200];
  assign t[161] = ~(t[200] | t[202]);
  assign t[162] = ~(x[7] | t[184]);
  assign t[163] = t[199] ? t[121] : t[122];
  assign t[164] = ~(t[79]);
  assign t[165] = t[199] ? t[124] : t[185];
  assign t[166] = ~(t[202] & t[162]);
  assign t[167] = ~(t[79] | t[199]);
  assign t[168] = ~(t[167] & t[186]);
  assign t[169] = ~(t[187] & t[188]);
  assign t[16] = ~(t[199] & t[200]);
  assign t[170] = ~(t[164] | t[189]);
  assign t[171] = t[199] ? t[166] : t[123];
  assign t[172] = ~(t[164] | t[190]);
  assign t[173] = ~(t[181] | t[177]);
  assign t[174] = ~(t[237]);
  assign t[175] = ~(t[232] | t[233]);
  assign t[176] = ~(t[164] | t[191]);
  assign t[177] = ~(t[164] | t[192]);
  assign t[178] = ~(t[31]);
  assign t[179] = ~(t[238]);
  assign t[17] = ~(t[201] & t[202]);
  assign t[180] = ~(t[235] | t[236]);
  assign t[181] = ~(t[164] | t[193]);
  assign t[182] = ~(t[194] & t[31]);
  assign t[183] = ~(t[164] | t[195]);
  assign t[184] = ~(t[200]);
  assign t[185] = ~(x[7] & t[187]);
  assign t[186] = ~(t[166] & t[185]);
  assign t[187] = ~(t[200] | t[159]);
  assign t[188] = t[164] & t[199];
  assign t[189] = t[199] ? t[196] : t[122];
  assign t[18] = x[7] ? t[27] : t[26];
  assign t[190] = t[199] ? t[197] : t[121];
  assign t[191] = t[199] ? t[123] : t[166];
  assign t[192] = t[199] ? t[122] : t[196];
  assign t[193] = t[199] ? t[185] : t[124];
  assign t[194] = ~(t[172] | t[51]);
  assign t[195] = t[199] ? t[121] : t[197];
  assign t[196] = ~(t[158] & t[202]);
  assign t[197] = ~(t[160] & t[202]);
  assign t[198] = (t[239]);
  assign t[199] = (t[240]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = ~(t[3]);
  assign t[200] = (t[241]);
  assign t[201] = (t[242]);
  assign t[202] = (t[243]);
  assign t[203] = (t[244]);
  assign t[204] = (t[245]);
  assign t[205] = (t[246]);
  assign t[206] = (t[247]);
  assign t[207] = (t[248]);
  assign t[208] = (t[249]);
  assign t[209] = (t[250]);
  assign t[20] = t[30] ? x[10] : x[9];
  assign t[210] = (t[251]);
  assign t[211] = (t[252]);
  assign t[212] = (t[253]);
  assign t[213] = (t[254]);
  assign t[214] = (t[255]);
  assign t[215] = (t[256]);
  assign t[216] = (t[257]);
  assign t[217] = (t[258]);
  assign t[218] = (t[259]);
  assign t[219] = (t[260]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[220] = (t[261]);
  assign t[221] = (t[262]);
  assign t[222] = (t[263]);
  assign t[223] = (t[264]);
  assign t[224] = (t[265]);
  assign t[225] = (t[266]);
  assign t[226] = (t[267]);
  assign t[227] = (t[268]);
  assign t[228] = (t[269]);
  assign t[229] = (t[270]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[230] = (t[271]);
  assign t[231] = (t[272]);
  assign t[232] = (t[273]);
  assign t[233] = (t[274]);
  assign t[234] = (t[275]);
  assign t[235] = (t[276]);
  assign t[236] = (t[277]);
  assign t[237] = (t[278]);
  assign t[238] = (t[279]);
  assign t[239] = t[280] ^ x[5];
  assign t[23] = ~(t[35] ^ t[36]);
  assign t[240] = t[281] ^ x[13];
  assign t[241] = t[282] ^ x[16];
  assign t[242] = t[283] ^ x[19];
  assign t[243] = t[284] ^ x[22];
  assign t[244] = t[285] ^ x[28];
  assign t[245] = t[286] ^ x[34];
  assign t[246] = t[287] ^ x[35];
  assign t[247] = t[288] ^ x[36];
  assign t[248] = t[289] ^ x[42];
  assign t[249] = t[290] ^ x[50];
  assign t[24] = x[7] ? t[38] : t[37];
  assign t[250] = t[291] ^ x[56];
  assign t[251] = t[292] ^ x[57];
  assign t[252] = t[293] ^ x[58];
  assign t[253] = t[294] ^ x[66];
  assign t[254] = t[295] ^ x[72];
  assign t[255] = t[296] ^ x[73];
  assign t[256] = t[297] ^ x[74];
  assign t[257] = t[298] ^ x[75];
  assign t[258] = t[299] ^ x[76];
  assign t[259] = t[300] ^ x[77];
  assign t[25] = x[7] ? t[40] : t[39];
  assign t[260] = t[301] ^ x[80];
  assign t[261] = t[302] ^ x[81];
  assign t[262] = t[303] ^ x[84];
  assign t[263] = t[304] ^ x[85];
  assign t[264] = t[305] ^ x[86];
  assign t[265] = t[306] ^ x[92];
  assign t[266] = t[307] ^ x[95];
  assign t[267] = t[308] ^ x[96];
  assign t[268] = t[309] ^ x[102];
  assign t[269] = t[310] ^ x[105];
  assign t[26] = ~(t[41] | t[42]);
  assign t[270] = t[311] ^ x[106];
  assign t[271] = t[312] ^ x[107];
  assign t[272] = t[313] ^ x[108];
  assign t[273] = t[314] ^ x[109];
  assign t[274] = t[315] ^ x[110];
  assign t[275] = t[316] ^ x[111];
  assign t[276] = t[317] ^ x[112];
  assign t[277] = t[318] ^ x[113];
  assign t[278] = t[319] ^ x[114];
  assign t[279] = t[320] ^ x[115];
  assign t[27] = ~(t[26] ^ t[43]);
  assign t[280] = (~t[321] & t[322]);
  assign t[281] = (~t[323] & t[324]);
  assign t[282] = (~t[325] & t[326]);
  assign t[283] = (~t[327] & t[328]);
  assign t[284] = (~t[329] & t[330]);
  assign t[285] = (~t[331] & t[332]);
  assign t[286] = (~t[333] & t[334]);
  assign t[287] = (~t[331] & t[335]);
  assign t[288] = (~t[331] & t[336]);
  assign t[289] = (~t[337] & t[338]);
  assign t[28] = x[7] ? t[45] : t[44];
  assign t[290] = (~t[339] & t[340]);
  assign t[291] = (~t[341] & t[342]);
  assign t[292] = (~t[333] & t[343]);
  assign t[293] = (~t[333] & t[344]);
  assign t[294] = (~t[345] & t[346]);
  assign t[295] = (~t[347] & t[348]);
  assign t[296] = (~t[331] & t[349]);
  assign t[297] = (~t[337] & t[350]);
  assign t[298] = (~t[337] & t[351]);
  assign t[299] = (~t[339] & t[352]);
  assign t[29] = x[7] ? t[47] : t[46];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (~t[339] & t[353]);
  assign t[301] = (~t[341] & t[354]);
  assign t[302] = (~t[341] & t[355]);
  assign t[303] = (~t[333] & t[356]);
  assign t[304] = (~t[345] & t[357]);
  assign t[305] = (~t[345] & t[358]);
  assign t[306] = (~t[359] & t[360]);
  assign t[307] = (~t[347] & t[361]);
  assign t[308] = (~t[347] & t[362]);
  assign t[309] = (~t[363] & t[364]);
  assign t[30] = ~(t[48]);
  assign t[310] = (~t[337] & t[365]);
  assign t[311] = (~t[339] & t[366]);
  assign t[312] = (~t[341] & t[367]);
  assign t[313] = (~t[345] & t[368]);
  assign t[314] = (~t[359] & t[369]);
  assign t[315] = (~t[359] & t[370]);
  assign t[316] = (~t[347] & t[371]);
  assign t[317] = (~t[363] & t[372]);
  assign t[318] = (~t[363] & t[373]);
  assign t[319] = (~t[359] & t[374]);
  assign t[31] = ~(t[49] | t[50]);
  assign t[320] = (~t[363] & t[375]);
  assign t[321] = t[376] ^ x[4];
  assign t[322] = t[377] ^ x[5];
  assign t[323] = t[378] ^ x[12];
  assign t[324] = t[379] ^ x[13];
  assign t[325] = t[380] ^ x[15];
  assign t[326] = t[381] ^ x[16];
  assign t[327] = t[382] ^ x[18];
  assign t[328] = t[383] ^ x[19];
  assign t[329] = t[384] ^ x[21];
  assign t[32] = ~(t[51] | t[52]);
  assign t[330] = t[385] ^ x[22];
  assign t[331] = t[386] ^ x[27];
  assign t[332] = t[387] ^ x[28];
  assign t[333] = t[388] ^ x[33];
  assign t[334] = t[389] ^ x[34];
  assign t[335] = t[390] ^ x[35];
  assign t[336] = t[391] ^ x[36];
  assign t[337] = t[392] ^ x[41];
  assign t[338] = t[393] ^ x[42];
  assign t[339] = t[394] ^ x[49];
  assign t[33] = ~(t[53] | t[54]);
  assign t[340] = t[395] ^ x[50];
  assign t[341] = t[396] ^ x[55];
  assign t[342] = t[397] ^ x[56];
  assign t[343] = t[398] ^ x[57];
  assign t[344] = t[399] ^ x[58];
  assign t[345] = t[400] ^ x[65];
  assign t[346] = t[401] ^ x[66];
  assign t[347] = t[402] ^ x[71];
  assign t[348] = t[403] ^ x[72];
  assign t[349] = t[404] ^ x[73];
  assign t[34] = ~(t[203] | t[55]);
  assign t[350] = t[405] ^ x[74];
  assign t[351] = t[406] ^ x[75];
  assign t[352] = t[407] ^ x[76];
  assign t[353] = t[408] ^ x[77];
  assign t[354] = t[409] ^ x[80];
  assign t[355] = t[410] ^ x[81];
  assign t[356] = t[411] ^ x[84];
  assign t[357] = t[412] ^ x[85];
  assign t[358] = t[413] ^ x[86];
  assign t[359] = t[414] ^ x[91];
  assign t[35] = ~(t[56] | t[57]);
  assign t[360] = t[415] ^ x[92];
  assign t[361] = t[416] ^ x[95];
  assign t[362] = t[417] ^ x[96];
  assign t[363] = t[418] ^ x[101];
  assign t[364] = t[419] ^ x[102];
  assign t[365] = t[420] ^ x[105];
  assign t[366] = t[421] ^ x[106];
  assign t[367] = t[422] ^ x[107];
  assign t[368] = t[423] ^ x[108];
  assign t[369] = t[424] ^ x[109];
  assign t[36] = ~(t[58] ^ t[59]);
  assign t[370] = t[425] ^ x[110];
  assign t[371] = t[426] ^ x[111];
  assign t[372] = t[427] ^ x[112];
  assign t[373] = t[428] ^ x[113];
  assign t[374] = t[429] ^ x[114];
  assign t[375] = t[430] ^ x[115];
  assign t[376] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[377] = (x[0]);
  assign t[378] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[379] = (x[11]);
  assign t[37] = ~(t[60] | t[61]);
  assign t[380] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[381] = (x[14]);
  assign t[382] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[383] = (x[17]);
  assign t[384] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[385] = (x[20]);
  assign t[386] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[387] = (x[24]);
  assign t[388] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[389] = (x[30]);
  assign t[38] = ~(t[39] ^ t[62]);
  assign t[390] = (x[25]);
  assign t[391] = (x[26]);
  assign t[392] = (x[37] & ~x[38] & ~x[39] & ~x[40]) | (~x[37] & x[38] & ~x[39] & ~x[40]) | (~x[37] & ~x[38] & x[39] & ~x[40]) | (~x[37] & ~x[38] & ~x[39] & x[40]) | (x[37] & x[38] & x[39] & ~x[40]) | (x[37] & x[38] & ~x[39] & x[40]) | (x[37] & ~x[38] & x[39] & x[40]) | (~x[37] & x[38] & x[39] & x[40]);
  assign t[393] = (x[38]);
  assign t[394] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[395] = (x[46]);
  assign t[396] = (x[51] & ~x[52] & ~x[53] & ~x[54]) | (~x[51] & x[52] & ~x[53] & ~x[54]) | (~x[51] & ~x[52] & x[53] & ~x[54]) | (~x[51] & ~x[52] & ~x[53] & x[54]) | (x[51] & x[52] & x[53] & ~x[54]) | (x[51] & x[52] & ~x[53] & x[54]) | (x[51] & ~x[52] & x[53] & x[54]) | (~x[51] & x[52] & x[53] & x[54]);
  assign t[397] = (x[52]);
  assign t[398] = (x[31]);
  assign t[399] = (x[32]);
  assign t[39] = ~(t[63] | t[64]);
  assign t[3] = ~(t[6]);
  assign t[400] = (x[61] & ~x[62] & ~x[63] & ~x[64]) | (~x[61] & x[62] & ~x[63] & ~x[64]) | (~x[61] & ~x[62] & x[63] & ~x[64]) | (~x[61] & ~x[62] & ~x[63] & x[64]) | (x[61] & x[62] & x[63] & ~x[64]) | (x[61] & x[62] & ~x[63] & x[64]) | (x[61] & ~x[62] & x[63] & x[64]) | (~x[61] & x[62] & x[63] & x[64]);
  assign t[401] = (x[62]);
  assign t[402] = (x[67] & ~x[68] & ~x[69] & ~x[70]) | (~x[67] & x[68] & ~x[69] & ~x[70]) | (~x[67] & ~x[68] & x[69] & ~x[70]) | (~x[67] & ~x[68] & ~x[69] & x[70]) | (x[67] & x[68] & x[69] & ~x[70]) | (x[67] & x[68] & ~x[69] & x[70]) | (x[67] & ~x[68] & x[69] & x[70]) | (~x[67] & x[68] & x[69] & x[70]);
  assign t[403] = (x[68]);
  assign t[404] = (x[23]);
  assign t[405] = (x[39]);
  assign t[406] = (x[40]);
  assign t[407] = (x[47]);
  assign t[408] = (x[48]);
  assign t[409] = (x[53]);
  assign t[40] = ~(t[44] ^ t[65]);
  assign t[410] = (x[54]);
  assign t[411] = (x[29]);
  assign t[412] = (x[63]);
  assign t[413] = (x[64]);
  assign t[414] = (x[87] & ~x[88] & ~x[89] & ~x[90]) | (~x[87] & x[88] & ~x[89] & ~x[90]) | (~x[87] & ~x[88] & x[89] & ~x[90]) | (~x[87] & ~x[88] & ~x[89] & x[90]) | (x[87] & x[88] & x[89] & ~x[90]) | (x[87] & x[88] & ~x[89] & x[90]) | (x[87] & ~x[88] & x[89] & x[90]) | (~x[87] & x[88] & x[89] & x[90]);
  assign t[415] = (x[88]);
  assign t[416] = (x[69]);
  assign t[417] = (x[70]);
  assign t[418] = (x[97] & ~x[98] & ~x[99] & ~x[100]) | (~x[97] & x[98] & ~x[99] & ~x[100]) | (~x[97] & ~x[98] & x[99] & ~x[100]) | (~x[97] & ~x[98] & ~x[99] & x[100]) | (x[97] & x[98] & x[99] & ~x[100]) | (x[97] & x[98] & ~x[99] & x[100]) | (x[97] & ~x[98] & x[99] & x[100]) | (~x[97] & x[98] & x[99] & x[100]);
  assign t[419] = (x[98]);
  assign t[41] = ~(t[66] | t[67]);
  assign t[420] = (x[37]);
  assign t[421] = (x[45]);
  assign t[422] = (x[51]);
  assign t[423] = (x[61]);
  assign t[424] = (x[89]);
  assign t[425] = (x[90]);
  assign t[426] = (x[67]);
  assign t[427] = (x[99]);
  assign t[428] = (x[100]);
  assign t[429] = (x[87]);
  assign t[42] = ~(t[204] | t[68]);
  assign t[430] = (x[97]);
  assign t[43] = ~(t[69] ^ t[70]);
  assign t[44] = ~(t[71] | t[72]);
  assign t[45] = ~(t[73] ^ t[74]);
  assign t[46] = ~(t[75] | t[76]);
  assign t[47] = ~(t[77] ^ t[78]);
  assign t[48] = ~(t[201]);
  assign t[49] = ~(t[79] | t[80]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[79] | t[81]);
  assign t[51] = ~(t[82] & t[83]);
  assign t[52] = ~(t[84] & t[85]);
  assign t[53] = ~(t[205]);
  assign t[54] = ~(t[206]);
  assign t[55] = ~(t[86] | t[87]);
  assign t[56] = ~(t[88] | t[89]);
  assign t[57] = ~(t[207] | t[90]);
  assign t[58] = t[91] ? x[44] : x[43];
  assign t[59] = ~(t[92] & t[84]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[93] | t[94]);
  assign t[61] = ~(t[208] | t[95]);
  assign t[62] = ~(t[96] ^ t[97]);
  assign t[63] = ~(t[98] | t[99]);
  assign t[64] = ~(t[209] | t[100]);
  assign t[65] = ~(t[101] ^ t[102]);
  assign t[66] = ~(t[210]);
  assign t[67] = ~(t[211]);
  assign t[68] = ~(t[103] | t[104]);
  assign t[69] = t[30] ? x[60] : x[59];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[105] & t[106]);
  assign t[71] = ~(t[107] | t[108]);
  assign t[72] = ~(t[212] | t[109]);
  assign t[73] = ~(t[110] | t[111]);
  assign t[74] = ~(t[112] ^ t[113]);
  assign t[75] = ~(t[114] | t[115]);
  assign t[76] = ~(t[213] | t[116]);
  assign t[77] = ~(t[117] | t[118]);
  assign t[78] = ~(t[119] ^ t[120]);
  assign t[79] = ~(t[201]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[199] ? t[122] : t[121];
  assign t[81] = t[199] ? t[124] : t[123];
  assign t[82] = ~(t[125] | t[126]);
  assign t[83] = ~(t[79] & t[127]);
  assign t[84] = ~(t[128] & t[129]);
  assign t[85] = t[79] | t[130];
  assign t[86] = ~(t[214]);
  assign t[87] = ~(t[205] | t[206]);
  assign t[88] = ~(t[215]);
  assign t[89] = ~(t[216]);
  assign t[8] = ~(t[14] ^ t[15]);
  assign t[90] = ~(t[131] | t[132]);
  assign t[91] = ~(t[48]);
  assign t[92] = ~(t[133] | t[134]);
  assign t[93] = ~(t[217]);
  assign t[94] = ~(t[218]);
  assign t[95] = ~(t[135] | t[136]);
  assign t[96] = t[137] ? x[79] : x[78];
  assign t[97] = t[138] | t[139];
  assign t[98] = ~(t[219]);
  assign t[99] = ~(t[220]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [112:0] x;
 output y;

 wire [446:0] t;
  assign t[0] = t[1] ? t[2] : t[265];
  assign t[100] = ~(t[289]);
  assign t[101] = ~(t[282] | t[283]);
  assign t[102] = ~(t[290]);
  assign t[103] = ~(t[291]);
  assign t[104] = ~(t[125] | t[126]);
  assign t[105] = ~(t[34]);
  assign t[106] = ~(t[85] | t[127]);
  assign t[107] = ~(t[128]);
  assign t[108] = x[7] & t[267];
  assign t[109] = ~(t[269]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = ~(x[7] | t[267]);
  assign t[111] = ~(t[267] | t[269]);
  assign t[112] = ~(x[7] | t[129]);
  assign t[113] = t[266] ? t[130] : t[84];
  assign t[114] = t[266] ? t[81] : t[131];
  assign t[115] = t[266] ? t[81] : t[82];
  assign t[116] = ~(t[35] | t[132]);
  assign t[117] = ~(t[54] & t[133]);
  assign t[118] = ~(t[123] & t[134]);
  assign t[119] = t[54] | t[135];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[292]);
  assign t[121] = ~(t[287] | t[288]);
  assign t[122] = ~(t[58] | t[136]);
  assign t[123] = t[269] & t[137];
  assign t[124] = ~(t[65]);
  assign t[125] = ~(t[293]);
  assign t[126] = ~(t[290] | t[291]);
  assign t[127] = ~(t[138] & t[65]);
  assign t[128] = ~(t[58] | t[139]);
  assign t[129] = ~(t[267]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[130] = ~(x[7] & t[140]);
  assign t[131] = ~(t[110] & t[269]);
  assign t[132] = ~(t[58] | t[141]);
  assign t[133] = ~(t[83] & t[87]);
  assign t[134] = t[110] | t[108];
  assign t[135] = t[266] ? t[83] : t[84];
  assign t[136] = t[266] ? t[83] : t[87];
  assign t[137] = ~(t[54] | t[266]);
  assign t[138] = ~(t[142] | t[91]);
  assign t[139] = t[266] ? t[82] : t[143];
  assign t[13] = x[7] ? t[20] : t[19];
  assign t[140] = ~(t[267] | t[109]);
  assign t[141] = t[266] ? t[84] : t[130];
  assign t[142] = ~(t[58] | t[144]);
  assign t[143] = ~(t[108] & t[269]);
  assign t[144] = t[266] ? t[143] : t[82];
  assign t[145] = t[1] ? t[146] : t[294];
  assign t[146] = x[6] ? t[148] : t[147];
  assign t[147] = x[7] ? t[150] : t[149];
  assign t[148] = t[151] ^ x[84];
  assign t[149] = t[152] ^ t[150];
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = ~(t[153] ^ t[154]);
  assign t[151] = x[85] ^ x[86];
  assign t[152] = t[23] ? x[86] : x[85];
  assign t[153] = x[7] ? t[156] : t[155];
  assign t[154] = ~(t[157] ^ t[158]);
  assign t[155] = ~(t[159] & t[160]);
  assign t[156] = t[161] ^ t[162];
  assign t[157] = x[7] ? t[164] : t[163];
  assign t[158] = x[7] ? t[166] : t[165];
  assign t[159] = ~(t[271] & t[40]);
  assign t[15] = ~(t[266] & t[267]);
  assign t[160] = ~(t[276] & t[167]);
  assign t[161] = t[23] ? x[88] : x[87];
  assign t[162] = ~(t[168] & t[169]);
  assign t[163] = ~(t[170] & t[171]);
  assign t[164] = t[172] ^ t[173];
  assign t[165] = ~(t[174] & t[175]);
  assign t[166] = t[176] ^ t[177];
  assign t[167] = ~(t[272] & t[39]);
  assign t[168] = ~(t[277] & t[63]);
  assign t[169] = ~(t[285] & t[178]);
  assign t[16] = ~(t[268] & t[269]);
  assign t[170] = ~(t[282] & t[75]);
  assign t[171] = ~(t[289] & t[179]);
  assign t[172] = t[105] ? x[90] : x[89];
  assign t[173] = ~(t[180] & t[181]);
  assign t[174] = ~(t[279] & t[68]);
  assign t[175] = ~(t[286] & t[182]);
  assign t[176] = t[23] ? x[92] : x[91];
  assign t[177] = ~(t[183] & t[184]);
  assign t[178] = ~(t[278] & t[62]);
  assign t[179] = ~(t[283] & t[74]);
  assign t[17] = t[23] ? x[10] : x[9];
  assign t[180] = ~(t[290] & t[103]);
  assign t[181] = ~(t[293] & t[185]);
  assign t[182] = ~(t[280] & t[67]);
  assign t[183] = ~(t[287] & t[96]);
  assign t[184] = ~(t[292] & t[186]);
  assign t[185] = ~(t[291] & t[102]);
  assign t[186] = ~(t[288] & t[95]);
  assign t[187] = t[1] ? t[188] : t[295];
  assign t[188] = x[6] ? t[190] : t[189];
  assign t[189] = x[7] ? t[192] : t[191];
  assign t[18] = ~(t[24] & t[25]);
  assign t[190] = t[193] ^ x[94];
  assign t[191] = t[194] ^ t[192];
  assign t[192] = ~(t[195] ^ t[196]);
  assign t[193] = x[95] ^ x[96];
  assign t[194] = t[23] ? x[96] : x[95];
  assign t[195] = x[7] ? t[198] : t[197];
  assign t[196] = ~(t[199] ^ t[200]);
  assign t[197] = ~(t[201] & t[202]);
  assign t[198] = t[203] ^ t[204];
  assign t[199] = x[7] ? t[206] : t[205];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = x[7] ? t[208] : t[207];
  assign t[201] = ~(t[40] & t[60]);
  assign t[202] = ~(t[209] & t[270]);
  assign t[203] = t[23] ? x[98] : x[97];
  assign t[204] = ~(t[210] & t[211]);
  assign t[205] = ~(t[212] & t[213]);
  assign t[206] = t[214] ^ t[215];
  assign t[207] = ~(t[216] & t[217]);
  assign t[208] = t[218] ^ t[219];
  assign t[209] = ~(t[220] & t[39]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = ~(t[63] & t[88]);
  assign t[211] = ~(t[221] & t[273]);
  assign t[212] = ~(t[75] & t[100]);
  assign t[213] = ~(t[222] & t[275]);
  assign t[214] = t[105] ? x[100] : x[99];
  assign t[215] = ~(t[223] & t[224]);
  assign t[216] = ~(t[68] & t[93]);
  assign t[217] = ~(t[225] & t[274]);
  assign t[218] = t[23] ? x[102] : x[101];
  assign t[219] = ~(t[226] & t[227]);
  assign t[21] = x[7] ? t[31] : t[30];
  assign t[220] = ~(t[276] & t[272]);
  assign t[221] = ~(t[228] & t[62]);
  assign t[222] = ~(t[229] & t[74]);
  assign t[223] = ~(t[103] & t[125]);
  assign t[224] = ~(t[230] & t[284]);
  assign t[225] = ~(t[231] & t[67]);
  assign t[226] = ~(t[96] & t[120]);
  assign t[227] = ~(t[232] & t[281]);
  assign t[228] = ~(t[285] & t[278]);
  assign t[229] = ~(t[289] & t[283]);
  assign t[22] = x[7] ? t[33] : t[32];
  assign t[230] = ~(t[233] & t[102]);
  assign t[231] = ~(t[286] & t[280]);
  assign t[232] = ~(t[234] & t[95]);
  assign t[233] = ~(t[293] & t[291]);
  assign t[234] = ~(t[292] & t[288]);
  assign t[235] = t[1] ? t[236] : t[296];
  assign t[236] = x[6] ? t[238] : t[237];
  assign t[237] = x[7] ? t[240] : t[239];
  assign t[238] = t[241] ^ x[104];
  assign t[239] = t[242] ^ t[240];
  assign t[23] = ~(t[34]);
  assign t[240] = ~(t[243] ^ t[244]);
  assign t[241] = x[105] ^ x[106];
  assign t[242] = t[23] ? x[106] : x[105];
  assign t[243] = x[7] ? t[246] : t[245];
  assign t[244] = ~(t[247] ^ t[248]);
  assign t[245] = ~(t[201] & t[249]);
  assign t[246] = t[250] ^ t[251];
  assign t[247] = x[7] ? t[253] : t[252];
  assign t[248] = x[7] ? t[255] : t[254];
  assign t[249] = t[26] | t[270];
  assign t[24] = ~(t[35] | t[36]);
  assign t[250] = t[23] ? x[108] : x[107];
  assign t[251] = ~(t[210] & t[256]);
  assign t[252] = ~(t[212] & t[257]);
  assign t[253] = t[258] ^ t[259];
  assign t[254] = ~(t[216] & t[260]);
  assign t[255] = t[261] ^ t[262];
  assign t[256] = t[42] | t[273];
  assign t[257] = t[50] | t[275];
  assign t[258] = t[105] ? x[110] : x[109];
  assign t[259] = ~(t[223] & t[263]);
  assign t[25] = ~(t[37] | t[38]);
  assign t[260] = t[46] | t[274];
  assign t[261] = t[23] ? x[112] : x[111];
  assign t[262] = ~(t[226] & t[264]);
  assign t[263] = t[77] | t[284];
  assign t[264] = t[70] | t[281];
  assign t[265] = (t[297]);
  assign t[266] = (t[298]);
  assign t[267] = (t[299]);
  assign t[268] = (t[300]);
  assign t[269] = (t[301]);
  assign t[26] = ~(t[39] | t[40]);
  assign t[270] = (t[302]);
  assign t[271] = (t[303]);
  assign t[272] = (t[304]);
  assign t[273] = (t[305]);
  assign t[274] = (t[306]);
  assign t[275] = (t[307]);
  assign t[276] = (t[308]);
  assign t[277] = (t[309]);
  assign t[278] = (t[310]);
  assign t[279] = (t[311]);
  assign t[27] = ~(t[270] | t[41]);
  assign t[280] = (t[312]);
  assign t[281] = (t[313]);
  assign t[282] = (t[314]);
  assign t[283] = (t[315]);
  assign t[284] = (t[316]);
  assign t[285] = (t[317]);
  assign t[286] = (t[318]);
  assign t[287] = (t[319]);
  assign t[288] = (t[320]);
  assign t[289] = (t[321]);
  assign t[28] = ~(t[42] | t[43]);
  assign t[290] = (t[322]);
  assign t[291] = (t[323]);
  assign t[292] = (t[324]);
  assign t[293] = (t[325]);
  assign t[294] = (t[326]);
  assign t[295] = (t[327]);
  assign t[296] = (t[328]);
  assign t[297] = t[329] ^ x[5];
  assign t[298] = t[330] ^ x[13];
  assign t[299] = t[331] ^ x[16];
  assign t[29] = ~(t[44] ^ t[45]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = t[332] ^ x[19];
  assign t[301] = t[333] ^ x[22];
  assign t[302] = t[334] ^ x[28];
  assign t[303] = t[335] ^ x[29];
  assign t[304] = t[336] ^ x[30];
  assign t[305] = t[337] ^ x[36];
  assign t[306] = t[338] ^ x[44];
  assign t[307] = t[339] ^ x[50];
  assign t[308] = t[340] ^ x[51];
  assign t[309] = t[341] ^ x[52];
  assign t[30] = ~(t[46] | t[47]);
  assign t[310] = t[342] ^ x[53];
  assign t[311] = t[343] ^ x[54];
  assign t[312] = t[344] ^ x[55];
  assign t[313] = t[345] ^ x[61];
  assign t[314] = t[346] ^ x[64];
  assign t[315] = t[347] ^ x[65];
  assign t[316] = t[348] ^ x[71];
  assign t[317] = t[349] ^ x[74];
  assign t[318] = t[350] ^ x[75];
  assign t[319] = t[351] ^ x[76];
  assign t[31] = ~(t[48] ^ t[49]);
  assign t[320] = t[352] ^ x[77];
  assign t[321] = t[353] ^ x[78];
  assign t[322] = t[354] ^ x[79];
  assign t[323] = t[355] ^ x[80];
  assign t[324] = t[356] ^ x[81];
  assign t[325] = t[357] ^ x[82];
  assign t[326] = t[358] ^ x[83];
  assign t[327] = t[359] ^ x[93];
  assign t[328] = t[360] ^ x[103];
  assign t[329] = (~t[361] & t[362]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[330] = (~t[363] & t[364]);
  assign t[331] = (~t[365] & t[366]);
  assign t[332] = (~t[367] & t[368]);
  assign t[333] = (~t[369] & t[370]);
  assign t[334] = (~t[371] & t[372]);
  assign t[335] = (~t[371] & t[373]);
  assign t[336] = (~t[371] & t[374]);
  assign t[337] = (~t[375] & t[376]);
  assign t[338] = (~t[377] & t[378]);
  assign t[339] = (~t[379] & t[380]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[340] = (~t[371] & t[381]);
  assign t[341] = (~t[375] & t[382]);
  assign t[342] = (~t[375] & t[383]);
  assign t[343] = (~t[377] & t[384]);
  assign t[344] = (~t[377] & t[385]);
  assign t[345] = (~t[386] & t[387]);
  assign t[346] = (~t[379] & t[388]);
  assign t[347] = (~t[379] & t[389]);
  assign t[348] = (~t[390] & t[391]);
  assign t[349] = (~t[375] & t[392]);
  assign t[34] = ~(t[268]);
  assign t[350] = (~t[377] & t[393]);
  assign t[351] = (~t[386] & t[394]);
  assign t[352] = (~t[386] & t[395]);
  assign t[353] = (~t[379] & t[396]);
  assign t[354] = (~t[390] & t[397]);
  assign t[355] = (~t[390] & t[398]);
  assign t[356] = (~t[386] & t[399]);
  assign t[357] = (~t[390] & t[400]);
  assign t[358] = (~t[361] & t[401]);
  assign t[359] = (~t[361] & t[402]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[360] = (~t[361] & t[403]);
  assign t[361] = t[404] ^ x[4];
  assign t[362] = t[405] ^ x[5];
  assign t[363] = t[406] ^ x[12];
  assign t[364] = t[407] ^ x[13];
  assign t[365] = t[408] ^ x[15];
  assign t[366] = t[409] ^ x[16];
  assign t[367] = t[410] ^ x[18];
  assign t[368] = t[411] ^ x[19];
  assign t[369] = t[412] ^ x[21];
  assign t[36] = ~(t[54] | t[56]);
  assign t[370] = t[413] ^ x[22];
  assign t[371] = t[414] ^ x[27];
  assign t[372] = t[415] ^ x[28];
  assign t[373] = t[416] ^ x[29];
  assign t[374] = t[417] ^ x[30];
  assign t[375] = t[418] ^ x[35];
  assign t[376] = t[419] ^ x[36];
  assign t[377] = t[420] ^ x[43];
  assign t[378] = t[421] ^ x[44];
  assign t[379] = t[422] ^ x[49];
  assign t[37] = ~(t[57]);
  assign t[380] = t[423] ^ x[50];
  assign t[381] = t[424] ^ x[51];
  assign t[382] = t[425] ^ x[52];
  assign t[383] = t[426] ^ x[53];
  assign t[384] = t[427] ^ x[54];
  assign t[385] = t[428] ^ x[55];
  assign t[386] = t[429] ^ x[60];
  assign t[387] = t[430] ^ x[61];
  assign t[388] = t[431] ^ x[64];
  assign t[389] = t[432] ^ x[65];
  assign t[38] = ~(t[58] | t[59]);
  assign t[390] = t[433] ^ x[70];
  assign t[391] = t[434] ^ x[71];
  assign t[392] = t[435] ^ x[74];
  assign t[393] = t[436] ^ x[75];
  assign t[394] = t[437] ^ x[76];
  assign t[395] = t[438] ^ x[77];
  assign t[396] = t[439] ^ x[78];
  assign t[397] = t[440] ^ x[79];
  assign t[398] = t[441] ^ x[80];
  assign t[399] = t[442] ^ x[81];
  assign t[39] = ~(t[271]);
  assign t[3] = ~(t[6]);
  assign t[400] = t[443] ^ x[82];
  assign t[401] = t[444] ^ x[83];
  assign t[402] = t[445] ^ x[93];
  assign t[403] = t[446] ^ x[103];
  assign t[404] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[405] = (x[0]);
  assign t[406] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[407] = (x[11]);
  assign t[408] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[409] = (x[14]);
  assign t[40] = ~(t[272]);
  assign t[410] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[411] = (x[17]);
  assign t[412] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[413] = (x[20]);
  assign t[414] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[415] = (x[24]);
  assign t[416] = (x[25]);
  assign t[417] = (x[26]);
  assign t[418] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[419] = (x[32]);
  assign t[41] = ~(t[60] | t[61]);
  assign t[420] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[421] = (x[40]);
  assign t[422] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[423] = (x[46]);
  assign t[424] = (x[23]);
  assign t[425] = (x[33]);
  assign t[426] = (x[34]);
  assign t[427] = (x[41]);
  assign t[428] = (x[42]);
  assign t[429] = (x[56] & ~x[57] & ~x[58] & ~x[59]) | (~x[56] & x[57] & ~x[58] & ~x[59]) | (~x[56] & ~x[57] & x[58] & ~x[59]) | (~x[56] & ~x[57] & ~x[58] & x[59]) | (x[56] & x[57] & x[58] & ~x[59]) | (x[56] & x[57] & ~x[58] & x[59]) | (x[56] & ~x[57] & x[58] & x[59]) | (~x[56] & x[57] & x[58] & x[59]);
  assign t[42] = ~(t[62] | t[63]);
  assign t[430] = (x[57]);
  assign t[431] = (x[47]);
  assign t[432] = (x[48]);
  assign t[433] = (x[66] & ~x[67] & ~x[68] & ~x[69]) | (~x[66] & x[67] & ~x[68] & ~x[69]) | (~x[66] & ~x[67] & x[68] & ~x[69]) | (~x[66] & ~x[67] & ~x[68] & x[69]) | (x[66] & x[67] & x[68] & ~x[69]) | (x[66] & x[67] & ~x[68] & x[69]) | (x[66] & ~x[67] & x[68] & x[69]) | (~x[66] & x[67] & x[68] & x[69]);
  assign t[434] = (x[67]);
  assign t[435] = (x[31]);
  assign t[436] = (x[39]);
  assign t[437] = (x[58]);
  assign t[438] = (x[59]);
  assign t[439] = (x[45]);
  assign t[43] = ~(t[273] | t[64]);
  assign t[440] = (x[68]);
  assign t[441] = (x[69]);
  assign t[442] = (x[56]);
  assign t[443] = (x[66]);
  assign t[444] = (x[1]);
  assign t[445] = (x[2]);
  assign t[446] = (x[3]);
  assign t[44] = t[23] ? x[38] : x[37];
  assign t[45] = ~(t[65] & t[66]);
  assign t[46] = ~(t[67] | t[68]);
  assign t[47] = ~(t[274] | t[69]);
  assign t[48] = ~(t[70] | t[71]);
  assign t[49] = ~(t[72] ^ t[73]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[74] | t[75]);
  assign t[51] = ~(t[275] | t[76]);
  assign t[52] = ~(t[77] | t[78]);
  assign t[53] = ~(t[79] ^ t[80]);
  assign t[54] = ~(t[268]);
  assign t[55] = t[266] ? t[82] : t[81];
  assign t[56] = t[266] ? t[84] : t[83];
  assign t[57] = ~(t[85] | t[86]);
  assign t[58] = ~(t[54]);
  assign t[59] = t[266] ? t[87] : t[83];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[276]);
  assign t[61] = ~(t[271] | t[272]);
  assign t[62] = ~(t[277]);
  assign t[63] = ~(t[278]);
  assign t[64] = ~(t[88] | t[89]);
  assign t[65] = ~(t[90] | t[36]);
  assign t[66] = ~(t[91] | t[92]);
  assign t[67] = ~(t[279]);
  assign t[68] = ~(t[280]);
  assign t[69] = ~(t[93] | t[94]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[95] | t[96]);
  assign t[71] = ~(t[281] | t[97]);
  assign t[72] = t[23] ? x[63] : x[62];
  assign t[73] = ~(t[98] & t[99]);
  assign t[74] = ~(t[282]);
  assign t[75] = ~(t[283]);
  assign t[76] = ~(t[100] | t[101]);
  assign t[77] = ~(t[102] | t[103]);
  assign t[78] = ~(t[284] | t[104]);
  assign t[79] = t[105] ? x[73] : x[72];
  assign t[7] = ~(t[8] ^ t[12]);
  assign t[80] = ~(t[106] & t[107]);
  assign t[81] = ~(t[108] & t[109]);
  assign t[82] = ~(t[110] & t[109]);
  assign t[83] = ~(x[7] & t[111]);
  assign t[84] = ~(t[112] & t[109]);
  assign t[85] = ~(t[58] | t[113]);
  assign t[86] = ~(t[58] | t[114]);
  assign t[87] = ~(t[269] & t[112]);
  assign t[88] = ~(t[285]);
  assign t[89] = ~(t[277] | t[278]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = ~(t[54] | t[115]);
  assign t[91] = ~(t[116] & t[117]);
  assign t[92] = ~(t[118] & t[119]);
  assign t[93] = ~(t[286]);
  assign t[94] = ~(t[279] | t[280]);
  assign t[95] = ~(t[287]);
  assign t[96] = ~(t[288]);
  assign t[97] = ~(t[120] | t[121]);
  assign t[98] = ~(t[122] | t[86]);
  assign t[99] = ~(t[123] | t[124]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0] & ~t[145] & ~t[187] & ~t[235]) | (~t[0] & t[145] & ~t[187] & ~t[235]) | (~t[0] & ~t[145] & t[187] & ~t[235]) | (~t[0] & ~t[145] & ~t[187] & t[235]) | (t[0] & t[145] & t[187] & ~t[235]) | (t[0] & t[145] & ~t[187] & t[235]) | (t[0] & ~t[145] & t[187] & t[235]) | (~t[0] & t[145] & t[187] & t[235]);
endmodule

module R2ind186(x, y);
 input [82:0] x;
 output y;

 wire [236:0] t;
  assign t[0] = t[1] ? t[2] : t[70];
  assign t[100] = t[129] ^ x[13];
  assign t[101] = t[130] ^ x[16];
  assign t[102] = t[131] ^ x[19];
  assign t[103] = t[132] ^ x[22];
  assign t[104] = t[133] ^ x[28];
  assign t[105] = t[134] ^ x[31];
  assign t[106] = t[135] ^ x[32];
  assign t[107] = t[136] ^ x[38];
  assign t[108] = t[137] ^ x[44];
  assign t[109] = t[138] ^ x[52];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[139] ^ x[55];
  assign t[111] = t[140] ^ x[56];
  assign t[112] = t[141] ^ x[57];
  assign t[113] = t[142] ^ x[58];
  assign t[114] = t[143] ^ x[59];
  assign t[115] = t[144] ^ x[65];
  assign t[116] = t[145] ^ x[66];
  assign t[117] = t[146] ^ x[67];
  assign t[118] = t[147] ^ x[73];
  assign t[119] = t[148] ^ x[74];
  assign t[11] = ~(x[6]);
  assign t[120] = t[149] ^ x[75];
  assign t[121] = t[150] ^ x[76];
  assign t[122] = t[151] ^ x[77];
  assign t[123] = t[152] ^ x[78];
  assign t[124] = t[153] ^ x[79];
  assign t[125] = t[154] ^ x[80];
  assign t[126] = t[155] ^ x[81];
  assign t[127] = t[156] ^ x[82];
  assign t[128] = (~t[157] & t[158]);
  assign t[129] = (~t[159] & t[160]);
  assign t[12] = t[17] ? x[10] : x[9];
  assign t[130] = (~t[161] & t[162]);
  assign t[131] = (~t[163] & t[164]);
  assign t[132] = (~t[165] & t[166]);
  assign t[133] = (~t[167] & t[168]);
  assign t[134] = (~t[167] & t[169]);
  assign t[135] = (~t[167] & t[170]);
  assign t[136] = (~t[171] & t[172]);
  assign t[137] = (~t[173] & t[174]);
  assign t[138] = (~t[175] & t[176]);
  assign t[139] = (~t[167] & t[177]);
  assign t[13] = x[7] ? t[19] : t[18];
  assign t[140] = (~t[171] & t[178]);
  assign t[141] = (~t[171] & t[179]);
  assign t[142] = (~t[173] & t[180]);
  assign t[143] = (~t[173] & t[181]);
  assign t[144] = (~t[182] & t[183]);
  assign t[145] = (~t[175] & t[184]);
  assign t[146] = (~t[175] & t[185]);
  assign t[147] = (~t[186] & t[187]);
  assign t[148] = (~t[171] & t[188]);
  assign t[149] = (~t[173] & t[189]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (~t[182] & t[190]);
  assign t[151] = (~t[182] & t[191]);
  assign t[152] = (~t[175] & t[192]);
  assign t[153] = (~t[186] & t[193]);
  assign t[154] = (~t[186] & t[194]);
  assign t[155] = (~t[182] & t[195]);
  assign t[156] = (~t[186] & t[196]);
  assign t[157] = t[197] ^ x[4];
  assign t[158] = t[198] ^ x[5];
  assign t[159] = t[199] ^ x[12];
  assign t[15] = ~(t[71] & t[72]);
  assign t[160] = t[200] ^ x[13];
  assign t[161] = t[201] ^ x[15];
  assign t[162] = t[202] ^ x[16];
  assign t[163] = t[203] ^ x[18];
  assign t[164] = t[204] ^ x[19];
  assign t[165] = t[205] ^ x[21];
  assign t[166] = t[206] ^ x[22];
  assign t[167] = t[207] ^ x[27];
  assign t[168] = t[208] ^ x[28];
  assign t[169] = t[209] ^ x[31];
  assign t[16] = ~(t[73] & t[74]);
  assign t[170] = t[210] ^ x[32];
  assign t[171] = t[211] ^ x[37];
  assign t[172] = t[212] ^ x[38];
  assign t[173] = t[213] ^ x[43];
  assign t[174] = t[214] ^ x[44];
  assign t[175] = t[215] ^ x[51];
  assign t[176] = t[216] ^ x[52];
  assign t[177] = t[217] ^ x[55];
  assign t[178] = t[218] ^ x[56];
  assign t[179] = t[219] ^ x[57];
  assign t[17] = ~(t[22]);
  assign t[180] = t[220] ^ x[58];
  assign t[181] = t[221] ^ x[59];
  assign t[182] = t[222] ^ x[64];
  assign t[183] = t[223] ^ x[65];
  assign t[184] = t[224] ^ x[66];
  assign t[185] = t[225] ^ x[67];
  assign t[186] = t[226] ^ x[72];
  assign t[187] = t[227] ^ x[73];
  assign t[188] = t[228] ^ x[74];
  assign t[189] = t[229] ^ x[75];
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = t[230] ^ x[76];
  assign t[191] = t[231] ^ x[77];
  assign t[192] = t[232] ^ x[78];
  assign t[193] = t[233] ^ x[79];
  assign t[194] = t[234] ^ x[80];
  assign t[195] = t[235] ^ x[81];
  assign t[196] = t[236] ^ x[82];
  assign t[197] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[198] = (x[3]);
  assign t[199] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (x[11]);
  assign t[201] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[202] = (x[14]);
  assign t[203] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[204] = (x[17]);
  assign t[205] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[206] = (x[20]);
  assign t[207] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[208] = (x[24]);
  assign t[209] = (x[26]);
  assign t[20] = x[7] ? t[28] : t[27];
  assign t[210] = (x[23]);
  assign t[211] = (x[33] & ~x[34] & ~x[35] & ~x[36]) | (~x[33] & x[34] & ~x[35] & ~x[36]) | (~x[33] & ~x[34] & x[35] & ~x[36]) | (~x[33] & ~x[34] & ~x[35] & x[36]) | (x[33] & x[34] & x[35] & ~x[36]) | (x[33] & x[34] & ~x[35] & x[36]) | (x[33] & ~x[34] & x[35] & x[36]) | (~x[33] & x[34] & x[35] & x[36]);
  assign t[212] = (x[34]);
  assign t[213] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[214] = (x[40]);
  assign t[215] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[216] = (x[48]);
  assign t[217] = (x[25]);
  assign t[218] = (x[36]);
  assign t[219] = (x[33]);
  assign t[21] = x[7] ? t[30] : t[29];
  assign t[220] = (x[42]);
  assign t[221] = (x[39]);
  assign t[222] = (x[60] & ~x[61] & ~x[62] & ~x[63]) | (~x[60] & x[61] & ~x[62] & ~x[63]) | (~x[60] & ~x[61] & x[62] & ~x[63]) | (~x[60] & ~x[61] & ~x[62] & x[63]) | (x[60] & x[61] & x[62] & ~x[63]) | (x[60] & x[61] & ~x[62] & x[63]) | (x[60] & ~x[61] & x[62] & x[63]) | (~x[60] & x[61] & x[62] & x[63]);
  assign t[223] = (x[61]);
  assign t[224] = (x[50]);
  assign t[225] = (x[47]);
  assign t[226] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[227] = (x[69]);
  assign t[228] = (x[35]);
  assign t[229] = (x[41]);
  assign t[22] = ~(t[73]);
  assign t[230] = (x[63]);
  assign t[231] = (x[60]);
  assign t[232] = (x[49]);
  assign t[233] = (x[71]);
  assign t[234] = (x[68]);
  assign t[235] = (x[62]);
  assign t[236] = (x[70]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = t[33] | t[75];
  assign t[25] = t[17] ? x[30] : x[29];
  assign t[26] = ~(t[34] & t[35]);
  assign t[27] = ~(t[36] & t[37]);
  assign t[28] = t[38] ^ t[39];
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[76]);
  assign t[32] = ~(t[77]);
  assign t[33] = ~(t[44] | t[31]);
  assign t[34] = ~(t[45] & t[46]);
  assign t[35] = t[47] | t[78];
  assign t[36] = ~(t[48] & t[49]);
  assign t[37] = t[50] | t[79];
  assign t[38] = t[51] ? x[46] : x[45];
  assign t[39] = ~(t[52] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[54] & t[55]);
  assign t[41] = t[56] | t[80];
  assign t[42] = t[17] ? x[54] : x[53];
  assign t[43] = ~(t[57] & t[58]);
  assign t[44] = ~(t[81]);
  assign t[45] = ~(t[82]);
  assign t[46] = ~(t[83]);
  assign t[47] = ~(t[59] | t[45]);
  assign t[48] = ~(t[84]);
  assign t[49] = ~(t[85]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[60] | t[48]);
  assign t[51] = ~(t[22]);
  assign t[52] = ~(t[61] & t[62]);
  assign t[53] = t[63] | t[86];
  assign t[54] = ~(t[87]);
  assign t[55] = ~(t[88]);
  assign t[56] = ~(t[64] | t[54]);
  assign t[57] = ~(t[65] & t[66]);
  assign t[58] = t[67] | t[89];
  assign t[59] = ~(t[90]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[91]);
  assign t[61] = ~(t[92]);
  assign t[62] = ~(t[93]);
  assign t[63] = ~(t[68] | t[61]);
  assign t[64] = ~(t[94]);
  assign t[65] = ~(t[95]);
  assign t[66] = ~(t[96]);
  assign t[67] = ~(t[69] | t[65]);
  assign t[68] = ~(t[97]);
  assign t[69] = ~(t[98]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[99]);
  assign t[71] = (t[100]);
  assign t[72] = (t[101]);
  assign t[73] = (t[102]);
  assign t[74] = (t[103]);
  assign t[75] = (t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = t[128] ^ x[5];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [82:0] x;
 output y;

 wire [242:0] t;
  assign t[0] = t[1] ? t[2] : t[76];
  assign t[100] = (t[129]);
  assign t[101] = (t[130]);
  assign t[102] = (t[131]);
  assign t[103] = (t[132]);
  assign t[104] = (t[133]);
  assign t[105] = t[134] ^ x[5];
  assign t[106] = t[135] ^ x[13];
  assign t[107] = t[136] ^ x[16];
  assign t[108] = t[137] ^ x[19];
  assign t[109] = t[138] ^ x[22];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[139] ^ x[28];
  assign t[111] = t[140] ^ x[31];
  assign t[112] = t[141] ^ x[32];
  assign t[113] = t[142] ^ x[38];
  assign t[114] = t[143] ^ x[44];
  assign t[115] = t[144] ^ x[52];
  assign t[116] = t[145] ^ x[55];
  assign t[117] = t[146] ^ x[56];
  assign t[118] = t[147] ^ x[57];
  assign t[119] = t[148] ^ x[58];
  assign t[11] = ~(x[6]);
  assign t[120] = t[149] ^ x[59];
  assign t[121] = t[150] ^ x[65];
  assign t[122] = t[151] ^ x[66];
  assign t[123] = t[152] ^ x[67];
  assign t[124] = t[153] ^ x[73];
  assign t[125] = t[154] ^ x[74];
  assign t[126] = t[155] ^ x[75];
  assign t[127] = t[156] ^ x[76];
  assign t[128] = t[157] ^ x[77];
  assign t[129] = t[158] ^ x[78];
  assign t[12] = t[17] ? x[10] : x[9];
  assign t[130] = t[159] ^ x[79];
  assign t[131] = t[160] ^ x[80];
  assign t[132] = t[161] ^ x[81];
  assign t[133] = t[162] ^ x[82];
  assign t[134] = (~t[163] & t[164]);
  assign t[135] = (~t[165] & t[166]);
  assign t[136] = (~t[167] & t[168]);
  assign t[137] = (~t[169] & t[170]);
  assign t[138] = (~t[171] & t[172]);
  assign t[139] = (~t[173] & t[174]);
  assign t[13] = x[7] ? t[19] : t[18];
  assign t[140] = (~t[173] & t[175]);
  assign t[141] = (~t[173] & t[176]);
  assign t[142] = (~t[177] & t[178]);
  assign t[143] = (~t[179] & t[180]);
  assign t[144] = (~t[181] & t[182]);
  assign t[145] = (~t[173] & t[183]);
  assign t[146] = (~t[177] & t[184]);
  assign t[147] = (~t[177] & t[185]);
  assign t[148] = (~t[179] & t[186]);
  assign t[149] = (~t[179] & t[187]);
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = (~t[188] & t[189]);
  assign t[151] = (~t[181] & t[190]);
  assign t[152] = (~t[181] & t[191]);
  assign t[153] = (~t[192] & t[193]);
  assign t[154] = (~t[177] & t[194]);
  assign t[155] = (~t[179] & t[195]);
  assign t[156] = (~t[188] & t[196]);
  assign t[157] = (~t[188] & t[197]);
  assign t[158] = (~t[181] & t[198]);
  assign t[159] = (~t[192] & t[199]);
  assign t[15] = ~(t[77] & t[78]);
  assign t[160] = (~t[192] & t[200]);
  assign t[161] = (~t[188] & t[201]);
  assign t[162] = (~t[192] & t[202]);
  assign t[163] = t[203] ^ x[4];
  assign t[164] = t[204] ^ x[5];
  assign t[165] = t[205] ^ x[12];
  assign t[166] = t[206] ^ x[13];
  assign t[167] = t[207] ^ x[15];
  assign t[168] = t[208] ^ x[16];
  assign t[169] = t[209] ^ x[18];
  assign t[16] = ~(t[79] & t[80]);
  assign t[170] = t[210] ^ x[19];
  assign t[171] = t[211] ^ x[21];
  assign t[172] = t[212] ^ x[22];
  assign t[173] = t[213] ^ x[27];
  assign t[174] = t[214] ^ x[28];
  assign t[175] = t[215] ^ x[31];
  assign t[176] = t[216] ^ x[32];
  assign t[177] = t[217] ^ x[37];
  assign t[178] = t[218] ^ x[38];
  assign t[179] = t[219] ^ x[43];
  assign t[17] = ~(t[22]);
  assign t[180] = t[220] ^ x[44];
  assign t[181] = t[221] ^ x[51];
  assign t[182] = t[222] ^ x[52];
  assign t[183] = t[223] ^ x[55];
  assign t[184] = t[224] ^ x[56];
  assign t[185] = t[225] ^ x[57];
  assign t[186] = t[226] ^ x[58];
  assign t[187] = t[227] ^ x[59];
  assign t[188] = t[228] ^ x[64];
  assign t[189] = t[229] ^ x[65];
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = t[230] ^ x[66];
  assign t[191] = t[231] ^ x[67];
  assign t[192] = t[232] ^ x[72];
  assign t[193] = t[233] ^ x[73];
  assign t[194] = t[234] ^ x[74];
  assign t[195] = t[235] ^ x[75];
  assign t[196] = t[236] ^ x[76];
  assign t[197] = t[237] ^ x[77];
  assign t[198] = t[238] ^ x[78];
  assign t[199] = t[239] ^ x[79];
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[80];
  assign t[201] = t[241] ^ x[81];
  assign t[202] = t[242] ^ x[82];
  assign t[203] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[204] = (x[2]);
  assign t[205] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[206] = (x[11]);
  assign t[207] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[208] = (x[14]);
  assign t[209] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[20] = x[7] ? t[28] : t[27];
  assign t[210] = (x[17]);
  assign t[211] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[212] = (x[20]);
  assign t[213] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[214] = (x[24]);
  assign t[215] = (x[26]);
  assign t[216] = (x[23]);
  assign t[217] = (x[33] & ~x[34] & ~x[35] & ~x[36]) | (~x[33] & x[34] & ~x[35] & ~x[36]) | (~x[33] & ~x[34] & x[35] & ~x[36]) | (~x[33] & ~x[34] & ~x[35] & x[36]) | (x[33] & x[34] & x[35] & ~x[36]) | (x[33] & x[34] & ~x[35] & x[36]) | (x[33] & ~x[34] & x[35] & x[36]) | (~x[33] & x[34] & x[35] & x[36]);
  assign t[218] = (x[34]);
  assign t[219] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[21] = x[7] ? t[30] : t[29];
  assign t[220] = (x[40]);
  assign t[221] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[222] = (x[48]);
  assign t[223] = (x[25]);
  assign t[224] = (x[36]);
  assign t[225] = (x[33]);
  assign t[226] = (x[42]);
  assign t[227] = (x[39]);
  assign t[228] = (x[60] & ~x[61] & ~x[62] & ~x[63]) | (~x[60] & x[61] & ~x[62] & ~x[63]) | (~x[60] & ~x[61] & x[62] & ~x[63]) | (~x[60] & ~x[61] & ~x[62] & x[63]) | (x[60] & x[61] & x[62] & ~x[63]) | (x[60] & x[61] & ~x[62] & x[63]) | (x[60] & ~x[61] & x[62] & x[63]) | (~x[60] & x[61] & x[62] & x[63]);
  assign t[229] = (x[61]);
  assign t[22] = ~(t[79]);
  assign t[230] = (x[50]);
  assign t[231] = (x[47]);
  assign t[232] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[233] = (x[69]);
  assign t[234] = (x[35]);
  assign t[235] = (x[41]);
  assign t[236] = (x[63]);
  assign t[237] = (x[60]);
  assign t[238] = (x[49]);
  assign t[239] = (x[71]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[240] = (x[68]);
  assign t[241] = (x[62]);
  assign t[242] = (x[70]);
  assign t[24] = ~(t[33] & t[81]);
  assign t[25] = t[17] ? x[30] : x[29];
  assign t[26] = ~(t[34] & t[35]);
  assign t[27] = ~(t[36] & t[37]);
  assign t[28] = t[38] ^ t[39];
  assign t[29] = ~(t[40] & t[41]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[82]);
  assign t[32] = ~(t[83]);
  assign t[33] = ~(t[44] & t[45]);
  assign t[34] = ~(t[46] & t[47]);
  assign t[35] = ~(t[48] & t[84]);
  assign t[36] = ~(t[49] & t[50]);
  assign t[37] = ~(t[51] & t[85]);
  assign t[38] = t[52] ? x[46] : x[45];
  assign t[39] = ~(t[53] & t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[55] & t[56]);
  assign t[41] = ~(t[57] & t[86]);
  assign t[42] = t[17] ? x[54] : x[53];
  assign t[43] = ~(t[58] & t[59]);
  assign t[44] = ~(t[83] & t[82]);
  assign t[45] = ~(t[87]);
  assign t[46] = ~(t[88]);
  assign t[47] = ~(t[89]);
  assign t[48] = ~(t[60] & t[61]);
  assign t[49] = ~(t[90]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[91]);
  assign t[51] = ~(t[62] & t[63]);
  assign t[52] = ~(t[22]);
  assign t[53] = ~(t[64] & t[65]);
  assign t[54] = ~(t[66] & t[92]);
  assign t[55] = ~(t[93]);
  assign t[56] = ~(t[94]);
  assign t[57] = ~(t[67] & t[68]);
  assign t[58] = ~(t[69] & t[70]);
  assign t[59] = ~(t[71] & t[95]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[89] & t[88]);
  assign t[61] = ~(t[96]);
  assign t[62] = ~(t[91] & t[90]);
  assign t[63] = ~(t[97]);
  assign t[64] = ~(t[98]);
  assign t[65] = ~(t[99]);
  assign t[66] = ~(t[72] & t[73]);
  assign t[67] = ~(t[94] & t[93]);
  assign t[68] = ~(t[100]);
  assign t[69] = ~(t[101]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[102]);
  assign t[71] = ~(t[74] & t[75]);
  assign t[72] = ~(t[99] & t[98]);
  assign t[73] = ~(t[103]);
  assign t[74] = ~(t[102] & t[101]);
  assign t[75] = ~(t[104]);
  assign t[76] = (t[105]);
  assign t[77] = (t[106]);
  assign t[78] = (t[107]);
  assign t[79] = (t[108]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[109]);
  assign t[81] = (t[110]);
  assign t[82] = (t[111]);
  assign t[83] = (t[112]);
  assign t[84] = (t[113]);
  assign t[85] = (t[114]);
  assign t[86] = (t[115]);
  assign t[87] = (t[116]);
  assign t[88] = (t[117]);
  assign t[89] = (t[118]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = (t[119]);
  assign t[91] = (t[120]);
  assign t[92] = (t[121]);
  assign t[93] = (t[122]);
  assign t[94] = (t[123]);
  assign t[95] = (t[124]);
  assign t[96] = (t[125]);
  assign t[97] = (t[126]);
  assign t[98] = (t[127]);
  assign t[99] = (t[128]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [76:0] x;
 output y;

 wire [200:0] t;
  assign t[0] = t[1] ? t[2] : t[64];
  assign t[100] = t[123] ^ x[55];
  assign t[101] = t[124] ^ x[58];
  assign t[102] = t[125] ^ x[59];
  assign t[103] = t[126] ^ x[65];
  assign t[104] = t[127] ^ x[66];
  assign t[105] = t[128] ^ x[67];
  assign t[106] = t[129] ^ x[73];
  assign t[107] = t[130] ^ x[74];
  assign t[108] = t[131] ^ x[75];
  assign t[109] = t[132] ^ x[76];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (~t[133] & t[134]);
  assign t[111] = (~t[135] & t[136]);
  assign t[112] = (~t[137] & t[138]);
  assign t[113] = (~t[139] & t[140]);
  assign t[114] = (~t[141] & t[142]);
  assign t[115] = (~t[143] & t[144]);
  assign t[116] = (~t[143] & t[145]);
  assign t[117] = (~t[143] & t[146]);
  assign t[118] = (~t[147] & t[148]);
  assign t[119] = (~t[147] & t[149]);
  assign t[11] = ~(x[6]);
  assign t[120] = (~t[150] & t[151]);
  assign t[121] = (~t[150] & t[152]);
  assign t[122] = (~t[153] & t[154]);
  assign t[123] = (~t[153] & t[155]);
  assign t[124] = (~t[147] & t[156]);
  assign t[125] = (~t[150] & t[157]);
  assign t[126] = (~t[158] & t[159]);
  assign t[127] = (~t[158] & t[160]);
  assign t[128] = (~t[153] & t[161]);
  assign t[129] = (~t[162] & t[163]);
  assign t[12] = t[17] ? x[10] : x[9];
  assign t[130] = (~t[162] & t[164]);
  assign t[131] = (~t[158] & t[165]);
  assign t[132] = (~t[162] & t[166]);
  assign t[133] = t[167] ^ x[4];
  assign t[134] = t[168] ^ x[5];
  assign t[135] = t[169] ^ x[12];
  assign t[136] = t[170] ^ x[13];
  assign t[137] = t[171] ^ x[15];
  assign t[138] = t[172] ^ x[16];
  assign t[139] = t[173] ^ x[18];
  assign t[13] = x[7] ? t[19] : t[18];
  assign t[140] = t[174] ^ x[19];
  assign t[141] = t[175] ^ x[21];
  assign t[142] = t[176] ^ x[22];
  assign t[143] = t[177] ^ x[27];
  assign t[144] = t[178] ^ x[28];
  assign t[145] = t[179] ^ x[29];
  assign t[146] = t[180] ^ x[32];
  assign t[147] = t[181] ^ x[37];
  assign t[148] = t[182] ^ x[38];
  assign t[149] = t[183] ^ x[39];
  assign t[14] = ~(t[20] ^ t[21]);
  assign t[150] = t[184] ^ x[44];
  assign t[151] = t[185] ^ x[45];
  assign t[152] = t[186] ^ x[46];
  assign t[153] = t[187] ^ x[53];
  assign t[154] = t[188] ^ x[54];
  assign t[155] = t[189] ^ x[55];
  assign t[156] = t[190] ^ x[58];
  assign t[157] = t[191] ^ x[59];
  assign t[158] = t[192] ^ x[64];
  assign t[159] = t[193] ^ x[65];
  assign t[15] = ~(t[65] & t[66]);
  assign t[160] = t[194] ^ x[66];
  assign t[161] = t[195] ^ x[67];
  assign t[162] = t[196] ^ x[72];
  assign t[163] = t[197] ^ x[73];
  assign t[164] = t[198] ^ x[74];
  assign t[165] = t[199] ^ x[75];
  assign t[166] = t[200] ^ x[76];
  assign t[167] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[168] = (x[1]);
  assign t[169] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[16] = ~(t[67] & t[68]);
  assign t[170] = (x[11]);
  assign t[171] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[172] = (x[14]);
  assign t[173] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[174] = (x[17]);
  assign t[175] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[176] = (x[20]);
  assign t[177] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[178] = (x[25]);
  assign t[179] = (x[23]);
  assign t[17] = ~(t[22]);
  assign t[180] = (x[26]);
  assign t[181] = (x[33] & ~x[34] & ~x[35] & ~x[36]) | (~x[33] & x[34] & ~x[35] & ~x[36]) | (~x[33] & ~x[34] & x[35] & ~x[36]) | (~x[33] & ~x[34] & ~x[35] & x[36]) | (x[33] & x[34] & x[35] & ~x[36]) | (x[33] & x[34] & ~x[35] & x[36]) | (x[33] & ~x[34] & x[35] & x[36]) | (~x[33] & x[34] & x[35] & x[36]);
  assign t[182] = (x[35]);
  assign t[183] = (x[33]);
  assign t[184] = (x[40] & ~x[41] & ~x[42] & ~x[43]) | (~x[40] & x[41] & ~x[42] & ~x[43]) | (~x[40] & ~x[41] & x[42] & ~x[43]) | (~x[40] & ~x[41] & ~x[42] & x[43]) | (x[40] & x[41] & x[42] & ~x[43]) | (x[40] & x[41] & ~x[42] & x[43]) | (x[40] & ~x[41] & x[42] & x[43]) | (~x[40] & x[41] & x[42] & x[43]);
  assign t[185] = (x[42]);
  assign t[186] = (x[40]);
  assign t[187] = (x[49] & ~x[50] & ~x[51] & ~x[52]) | (~x[49] & x[50] & ~x[51] & ~x[52]) | (~x[49] & ~x[50] & x[51] & ~x[52]) | (~x[49] & ~x[50] & ~x[51] & x[52]) | (x[49] & x[50] & x[51] & ~x[52]) | (x[49] & x[50] & ~x[51] & x[52]) | (x[49] & ~x[50] & x[51] & x[52]) | (~x[49] & x[50] & x[51] & x[52]);
  assign t[188] = (x[51]);
  assign t[189] = (x[49]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[190] = (x[36]);
  assign t[191] = (x[43]);
  assign t[192] = (x[60] & ~x[61] & ~x[62] & ~x[63]) | (~x[60] & x[61] & ~x[62] & ~x[63]) | (~x[60] & ~x[61] & x[62] & ~x[63]) | (~x[60] & ~x[61] & ~x[62] & x[63]) | (x[60] & x[61] & x[62] & ~x[63]) | (x[60] & x[61] & ~x[62] & x[63]) | (x[60] & ~x[61] & x[62] & x[63]) | (~x[60] & x[61] & x[62] & x[63]);
  assign t[193] = (x[62]);
  assign t[194] = (x[60]);
  assign t[195] = (x[52]);
  assign t[196] = (x[68] & ~x[69] & ~x[70] & ~x[71]) | (~x[68] & x[69] & ~x[70] & ~x[71]) | (~x[68] & ~x[69] & x[70] & ~x[71]) | (~x[68] & ~x[69] & ~x[70] & x[71]) | (x[68] & x[69] & x[70] & ~x[71]) | (x[68] & x[69] & ~x[70] & x[71]) | (x[68] & ~x[69] & x[70] & x[71]) | (~x[68] & x[69] & x[70] & x[71]);
  assign t[197] = (x[70]);
  assign t[198] = (x[68]);
  assign t[199] = (x[63]);
  assign t[19] = t[25] ^ t[26];
  assign t[1] = ~(t[3]);
  assign t[200] = (x[71]);
  assign t[20] = x[7] ? t[28] : t[27];
  assign t[21] = x[7] ? t[30] : t[29];
  assign t[22] = ~(t[67]);
  assign t[23] = ~(t[69] & t[31]);
  assign t[24] = ~(t[70] & t[32]);
  assign t[25] = t[17] ? x[31] : x[30];
  assign t[26] = ~(t[33] & t[34]);
  assign t[27] = ~(t[35] & t[36]);
  assign t[28] = t[37] ^ t[38];
  assign t[29] = ~(t[39] & t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[41] ^ t[42];
  assign t[31] = ~(t[71]);
  assign t[32] = ~(t[71] & t[43]);
  assign t[33] = ~(t[72] & t[44]);
  assign t[34] = ~(t[73] & t[45]);
  assign t[35] = ~(t[74] & t[46]);
  assign t[36] = ~(t[75] & t[47]);
  assign t[37] = t[48] ? x[48] : x[47];
  assign t[38] = ~(t[49] & t[50]);
  assign t[39] = ~(t[76] & t[51]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[77] & t[52]);
  assign t[41] = t[17] ? x[57] : x[56];
  assign t[42] = ~(t[53] & t[54]);
  assign t[43] = ~(t[69]);
  assign t[44] = ~(t[78]);
  assign t[45] = ~(t[78] & t[55]);
  assign t[46] = ~(t[79]);
  assign t[47] = ~(t[79] & t[56]);
  assign t[48] = ~(t[22]);
  assign t[49] = ~(t[80] & t[57]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[81] & t[58]);
  assign t[51] = ~(t[82]);
  assign t[52] = ~(t[82] & t[59]);
  assign t[53] = ~(t[83] & t[60]);
  assign t[54] = ~(t[84] & t[61]);
  assign t[55] = ~(t[72]);
  assign t[56] = ~(t[74]);
  assign t[57] = ~(t[85]);
  assign t[58] = ~(t[85] & t[62]);
  assign t[59] = ~(t[76]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[86]);
  assign t[61] = ~(t[86] & t[63]);
  assign t[62] = ~(t[80]);
  assign t[63] = ~(t[83]);
  assign t[64] = (t[87]);
  assign t[65] = (t[88]);
  assign t[66] = (t[89]);
  assign t[67] = (t[90]);
  assign t[68] = (t[91]);
  assign t[69] = (t[92]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[93]);
  assign t[71] = (t[94]);
  assign t[72] = (t[95]);
  assign t[73] = (t[96]);
  assign t[74] = (t[97]);
  assign t[75] = (t[98]);
  assign t[76] = (t[99]);
  assign t[77] = (t[100]);
  assign t[78] = (t[101]);
  assign t[79] = (t[102]);
  assign t[7] = t[12] ^ t[8];
  assign t[80] = (t[103]);
  assign t[81] = (t[104]);
  assign t[82] = (t[105]);
  assign t[83] = (t[106]);
  assign t[84] = (t[107]);
  assign t[85] = (t[108]);
  assign t[86] = (t[109]);
  assign t[87] = t[110] ^ x[5];
  assign t[88] = t[111] ^ x[13];
  assign t[89] = t[112] ^ x[16];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = t[113] ^ x[19];
  assign t[91] = t[114] ^ x[22];
  assign t[92] = t[115] ^ x[28];
  assign t[93] = t[116] ^ x[29];
  assign t[94] = t[117] ^ x[32];
  assign t[95] = t[118] ^ x[38];
  assign t[96] = t[119] ^ x[39];
  assign t[97] = t[120] ^ x[45];
  assign t[98] = t[121] ^ x[46];
  assign t[99] = t[122] ^ x[54];
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [82:0] x;
 output y;

 wire [311:0] t;
  assign t[0] = t[1] ? t[2] : t[145];
  assign t[100] = ~(t[169]);
  assign t[101] = ~(t[162] | t[163]);
  assign t[102] = ~(t[170]);
  assign t[103] = ~(t[171]);
  assign t[104] = ~(t[125] | t[126]);
  assign t[105] = ~(t[34]);
  assign t[106] = ~(t[85] | t[127]);
  assign t[107] = ~(t[128]);
  assign t[108] = x[7] & t[147];
  assign t[109] = ~(t[149]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = ~(x[7] | t[147]);
  assign t[111] = ~(t[147] | t[149]);
  assign t[112] = ~(x[7] | t[129]);
  assign t[113] = t[146] ? t[130] : t[84];
  assign t[114] = t[146] ? t[81] : t[131];
  assign t[115] = t[146] ? t[81] : t[82];
  assign t[116] = ~(t[35] | t[132]);
  assign t[117] = ~(t[54] & t[133]);
  assign t[118] = ~(t[123] & t[134]);
  assign t[119] = t[54] | t[135];
  assign t[11] = ~(x[6]);
  assign t[120] = ~(t[172]);
  assign t[121] = ~(t[167] | t[168]);
  assign t[122] = ~(t[58] | t[136]);
  assign t[123] = t[149] & t[137];
  assign t[124] = ~(t[65]);
  assign t[125] = ~(t[173]);
  assign t[126] = ~(t[170] | t[171]);
  assign t[127] = ~(t[138] & t[65]);
  assign t[128] = ~(t[58] | t[139]);
  assign t[129] = ~(t[147]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[130] = ~(x[7] & t[140]);
  assign t[131] = ~(t[110] & t[149]);
  assign t[132] = ~(t[58] | t[141]);
  assign t[133] = ~(t[83] & t[87]);
  assign t[134] = t[110] | t[108];
  assign t[135] = t[146] ? t[83] : t[84];
  assign t[136] = t[146] ? t[83] : t[87];
  assign t[137] = ~(t[54] | t[146]);
  assign t[138] = ~(t[142] | t[91]);
  assign t[139] = t[146] ? t[82] : t[143];
  assign t[13] = x[7] ? t[20] : t[19];
  assign t[140] = ~(t[147] | t[109]);
  assign t[141] = t[146] ? t[84] : t[130];
  assign t[142] = ~(t[58] | t[144]);
  assign t[143] = ~(t[108] & t[149]);
  assign t[144] = t[146] ? t[143] : t[82];
  assign t[145] = (t[174]);
  assign t[146] = (t[175]);
  assign t[147] = (t[176]);
  assign t[148] = (t[177]);
  assign t[149] = (t[178]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[150] = (t[179]);
  assign t[151] = (t[180]);
  assign t[152] = (t[181]);
  assign t[153] = (t[182]);
  assign t[154] = (t[183]);
  assign t[155] = (t[184]);
  assign t[156] = (t[185]);
  assign t[157] = (t[186]);
  assign t[158] = (t[187]);
  assign t[159] = (t[188]);
  assign t[15] = ~(t[146] & t[147]);
  assign t[160] = (t[189]);
  assign t[161] = (t[190]);
  assign t[162] = (t[191]);
  assign t[163] = (t[192]);
  assign t[164] = (t[193]);
  assign t[165] = (t[194]);
  assign t[166] = (t[195]);
  assign t[167] = (t[196]);
  assign t[168] = (t[197]);
  assign t[169] = (t[198]);
  assign t[16] = ~(t[148] & t[149]);
  assign t[170] = (t[199]);
  assign t[171] = (t[200]);
  assign t[172] = (t[201]);
  assign t[173] = (t[202]);
  assign t[174] = t[203] ^ x[5];
  assign t[175] = t[204] ^ x[13];
  assign t[176] = t[205] ^ x[16];
  assign t[177] = t[206] ^ x[19];
  assign t[178] = t[207] ^ x[22];
  assign t[179] = t[208] ^ x[28];
  assign t[17] = t[23] ? x[10] : x[9];
  assign t[180] = t[209] ^ x[29];
  assign t[181] = t[210] ^ x[30];
  assign t[182] = t[211] ^ x[36];
  assign t[183] = t[212] ^ x[44];
  assign t[184] = t[213] ^ x[50];
  assign t[185] = t[214] ^ x[51];
  assign t[186] = t[215] ^ x[52];
  assign t[187] = t[216] ^ x[53];
  assign t[188] = t[217] ^ x[54];
  assign t[189] = t[218] ^ x[55];
  assign t[18] = ~(t[24] & t[25]);
  assign t[190] = t[219] ^ x[61];
  assign t[191] = t[220] ^ x[64];
  assign t[192] = t[221] ^ x[65];
  assign t[193] = t[222] ^ x[71];
  assign t[194] = t[223] ^ x[74];
  assign t[195] = t[224] ^ x[75];
  assign t[196] = t[225] ^ x[76];
  assign t[197] = t[226] ^ x[77];
  assign t[198] = t[227] ^ x[78];
  assign t[199] = t[228] ^ x[79];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[229] ^ x[80];
  assign t[201] = t[230] ^ x[81];
  assign t[202] = t[231] ^ x[82];
  assign t[203] = (~t[232] & t[233]);
  assign t[204] = (~t[234] & t[235]);
  assign t[205] = (~t[236] & t[237]);
  assign t[206] = (~t[238] & t[239]);
  assign t[207] = (~t[240] & t[241]);
  assign t[208] = (~t[242] & t[243]);
  assign t[209] = (~t[242] & t[244]);
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = (~t[242] & t[245]);
  assign t[211] = (~t[246] & t[247]);
  assign t[212] = (~t[248] & t[249]);
  assign t[213] = (~t[250] & t[251]);
  assign t[214] = (~t[242] & t[252]);
  assign t[215] = (~t[246] & t[253]);
  assign t[216] = (~t[246] & t[254]);
  assign t[217] = (~t[248] & t[255]);
  assign t[218] = (~t[248] & t[256]);
  assign t[219] = (~t[257] & t[258]);
  assign t[21] = x[7] ? t[31] : t[30];
  assign t[220] = (~t[250] & t[259]);
  assign t[221] = (~t[250] & t[260]);
  assign t[222] = (~t[261] & t[262]);
  assign t[223] = (~t[246] & t[263]);
  assign t[224] = (~t[248] & t[264]);
  assign t[225] = (~t[257] & t[265]);
  assign t[226] = (~t[257] & t[266]);
  assign t[227] = (~t[250] & t[267]);
  assign t[228] = (~t[261] & t[268]);
  assign t[229] = (~t[261] & t[269]);
  assign t[22] = x[7] ? t[33] : t[32];
  assign t[230] = (~t[257] & t[270]);
  assign t[231] = (~t[261] & t[271]);
  assign t[232] = t[272] ^ x[4];
  assign t[233] = t[273] ^ x[5];
  assign t[234] = t[274] ^ x[12];
  assign t[235] = t[275] ^ x[13];
  assign t[236] = t[276] ^ x[15];
  assign t[237] = t[277] ^ x[16];
  assign t[238] = t[278] ^ x[18];
  assign t[239] = t[279] ^ x[19];
  assign t[23] = ~(t[34]);
  assign t[240] = t[280] ^ x[21];
  assign t[241] = t[281] ^ x[22];
  assign t[242] = t[282] ^ x[27];
  assign t[243] = t[283] ^ x[28];
  assign t[244] = t[284] ^ x[29];
  assign t[245] = t[285] ^ x[30];
  assign t[246] = t[286] ^ x[35];
  assign t[247] = t[287] ^ x[36];
  assign t[248] = t[288] ^ x[43];
  assign t[249] = t[289] ^ x[44];
  assign t[24] = ~(t[35] | t[36]);
  assign t[250] = t[290] ^ x[49];
  assign t[251] = t[291] ^ x[50];
  assign t[252] = t[292] ^ x[51];
  assign t[253] = t[293] ^ x[52];
  assign t[254] = t[294] ^ x[53];
  assign t[255] = t[295] ^ x[54];
  assign t[256] = t[296] ^ x[55];
  assign t[257] = t[297] ^ x[60];
  assign t[258] = t[298] ^ x[61];
  assign t[259] = t[299] ^ x[64];
  assign t[25] = ~(t[37] | t[38]);
  assign t[260] = t[300] ^ x[65];
  assign t[261] = t[301] ^ x[70];
  assign t[262] = t[302] ^ x[71];
  assign t[263] = t[303] ^ x[74];
  assign t[264] = t[304] ^ x[75];
  assign t[265] = t[305] ^ x[76];
  assign t[266] = t[306] ^ x[77];
  assign t[267] = t[307] ^ x[78];
  assign t[268] = t[308] ^ x[79];
  assign t[269] = t[309] ^ x[80];
  assign t[26] = ~(t[39] | t[40]);
  assign t[270] = t[310] ^ x[81];
  assign t[271] = t[311] ^ x[82];
  assign t[272] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[273] = (x[0]);
  assign t[274] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[275] = (x[11]);
  assign t[276] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[277] = (x[14]);
  assign t[278] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[279] = (x[17]);
  assign t[27] = ~(t[150] | t[41]);
  assign t[280] = (x[20] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[20] & 1'b0 & ~1'b0 & ~1'b0) | (~x[20] & ~1'b0 & 1'b0 & ~1'b0) | (~x[20] & ~1'b0 & ~1'b0 & 1'b0) | (x[20] & 1'b0 & 1'b0 & ~1'b0) | (x[20] & 1'b0 & ~1'b0 & 1'b0) | (x[20] & ~1'b0 & 1'b0 & 1'b0) | (~x[20] & 1'b0 & 1'b0 & 1'b0);
  assign t[281] = (x[20]);
  assign t[282] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[283] = (x[24]);
  assign t[284] = (x[25]);
  assign t[285] = (x[26]);
  assign t[286] = (x[31] & ~x[32] & ~x[33] & ~x[34]) | (~x[31] & x[32] & ~x[33] & ~x[34]) | (~x[31] & ~x[32] & x[33] & ~x[34]) | (~x[31] & ~x[32] & ~x[33] & x[34]) | (x[31] & x[32] & x[33] & ~x[34]) | (x[31] & x[32] & ~x[33] & x[34]) | (x[31] & ~x[32] & x[33] & x[34]) | (~x[31] & x[32] & x[33] & x[34]);
  assign t[287] = (x[32]);
  assign t[288] = (x[39] & ~x[40] & ~x[41] & ~x[42]) | (~x[39] & x[40] & ~x[41] & ~x[42]) | (~x[39] & ~x[40] & x[41] & ~x[42]) | (~x[39] & ~x[40] & ~x[41] & x[42]) | (x[39] & x[40] & x[41] & ~x[42]) | (x[39] & x[40] & ~x[41] & x[42]) | (x[39] & ~x[40] & x[41] & x[42]) | (~x[39] & x[40] & x[41] & x[42]);
  assign t[289] = (x[40]);
  assign t[28] = ~(t[42] | t[43]);
  assign t[290] = (x[45] & ~x[46] & ~x[47] & ~x[48]) | (~x[45] & x[46] & ~x[47] & ~x[48]) | (~x[45] & ~x[46] & x[47] & ~x[48]) | (~x[45] & ~x[46] & ~x[47] & x[48]) | (x[45] & x[46] & x[47] & ~x[48]) | (x[45] & x[46] & ~x[47] & x[48]) | (x[45] & ~x[46] & x[47] & x[48]) | (~x[45] & x[46] & x[47] & x[48]);
  assign t[291] = (x[46]);
  assign t[292] = (x[23]);
  assign t[293] = (x[33]);
  assign t[294] = (x[34]);
  assign t[295] = (x[41]);
  assign t[296] = (x[42]);
  assign t[297] = (x[56] & ~x[57] & ~x[58] & ~x[59]) | (~x[56] & x[57] & ~x[58] & ~x[59]) | (~x[56] & ~x[57] & x[58] & ~x[59]) | (~x[56] & ~x[57] & ~x[58] & x[59]) | (x[56] & x[57] & x[58] & ~x[59]) | (x[56] & x[57] & ~x[58] & x[59]) | (x[56] & ~x[57] & x[58] & x[59]) | (~x[56] & x[57] & x[58] & x[59]);
  assign t[298] = (x[57]);
  assign t[299] = (x[47]);
  assign t[29] = ~(t[44] ^ t[45]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[300] = (x[48]);
  assign t[301] = (x[66] & ~x[67] & ~x[68] & ~x[69]) | (~x[66] & x[67] & ~x[68] & ~x[69]) | (~x[66] & ~x[67] & x[68] & ~x[69]) | (~x[66] & ~x[67] & ~x[68] & x[69]) | (x[66] & x[67] & x[68] & ~x[69]) | (x[66] & x[67] & ~x[68] & x[69]) | (x[66] & ~x[67] & x[68] & x[69]) | (~x[66] & x[67] & x[68] & x[69]);
  assign t[302] = (x[67]);
  assign t[303] = (x[31]);
  assign t[304] = (x[39]);
  assign t[305] = (x[58]);
  assign t[306] = (x[59]);
  assign t[307] = (x[45]);
  assign t[308] = (x[68]);
  assign t[309] = (x[69]);
  assign t[30] = ~(t[46] | t[47]);
  assign t[310] = (x[56]);
  assign t[311] = (x[66]);
  assign t[31] = ~(t[48] ^ t[49]);
  assign t[32] = ~(t[50] | t[51]);
  assign t[33] = ~(t[52] ^ t[53]);
  assign t[34] = ~(t[148]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[36] = ~(t[54] | t[56]);
  assign t[37] = ~(t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = ~(t[151]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[152]);
  assign t[41] = ~(t[60] | t[61]);
  assign t[42] = ~(t[62] | t[63]);
  assign t[43] = ~(t[153] | t[64]);
  assign t[44] = t[23] ? x[38] : x[37];
  assign t[45] = ~(t[65] & t[66]);
  assign t[46] = ~(t[67] | t[68]);
  assign t[47] = ~(t[154] | t[69]);
  assign t[48] = ~(t[70] | t[71]);
  assign t[49] = ~(t[72] ^ t[73]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[74] | t[75]);
  assign t[51] = ~(t[155] | t[76]);
  assign t[52] = ~(t[77] | t[78]);
  assign t[53] = ~(t[79] ^ t[80]);
  assign t[54] = ~(t[148]);
  assign t[55] = t[146] ? t[82] : t[81];
  assign t[56] = t[146] ? t[84] : t[83];
  assign t[57] = ~(t[85] | t[86]);
  assign t[58] = ~(t[54]);
  assign t[59] = t[146] ? t[87] : t[83];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[156]);
  assign t[61] = ~(t[151] | t[152]);
  assign t[62] = ~(t[157]);
  assign t[63] = ~(t[158]);
  assign t[64] = ~(t[88] | t[89]);
  assign t[65] = ~(t[90] | t[36]);
  assign t[66] = ~(t[91] | t[92]);
  assign t[67] = ~(t[159]);
  assign t[68] = ~(t[160]);
  assign t[69] = ~(t[93] | t[94]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[95] | t[96]);
  assign t[71] = ~(t[161] | t[97]);
  assign t[72] = t[23] ? x[63] : x[62];
  assign t[73] = ~(t[98] & t[99]);
  assign t[74] = ~(t[162]);
  assign t[75] = ~(t[163]);
  assign t[76] = ~(t[100] | t[101]);
  assign t[77] = ~(t[102] | t[103]);
  assign t[78] = ~(t[164] | t[104]);
  assign t[79] = t[105] ? x[73] : x[72];
  assign t[7] = ~(t[8] ^ t[12]);
  assign t[80] = ~(t[106] & t[107]);
  assign t[81] = ~(t[108] & t[109]);
  assign t[82] = ~(t[110] & t[109]);
  assign t[83] = ~(x[7] & t[111]);
  assign t[84] = ~(t[112] & t[109]);
  assign t[85] = ~(t[58] | t[113]);
  assign t[86] = ~(t[58] | t[114]);
  assign t[87] = ~(t[149] & t[112]);
  assign t[88] = ~(t[165]);
  assign t[89] = ~(t[157] | t[158]);
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = ~(t[54] | t[115]);
  assign t[91] = ~(t[116] & t[117]);
  assign t[92] = ~(t[118] & t[119]);
  assign t[93] = ~(t[166]);
  assign t[94] = ~(t[159] | t[160]);
  assign t[95] = ~(t[167]);
  assign t[96] = ~(t[168]);
  assign t[97] = ~(t[120] | t[121]);
  assign t[98] = ~(t[122] | t[86]);
  assign t[99] = ~(t[123] | t[124]);
  assign t[9] = x[9] ^ x[10];
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [355:0] x;
 output [189:0] y;

  R2ind0 R2ind0_inst(.x({x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[5], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[5], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[5], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[5], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[5]));
  R2ind6 R2ind6_inst(.y(y[6]));
  R2ind7 R2ind7_inst(.y(y[7]));
  R2ind8 R2ind8_inst(.y(y[8]));
  R2ind9 R2ind9_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[11], x[10], x[9], x[18]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[11], x[10], x[9], x[18]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[11], x[10], x[9], x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[18]}), .y(y[15]));
  R2ind16 R2ind16_inst(.y(y[16]));
  R2ind17 R2ind17_inst(.y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.x({x[11], x[10], x[9], x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[18]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[18]}), .y(y[20]));
  R2ind21 R2ind21_inst(.y(y[21]));
  R2ind22 R2ind22_inst(.y(y[22]));
  R2ind23 R2ind23_inst(.y(y[23]));
  R2ind24 R2ind24_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[18]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[18]}), .y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.y(y[28]));
  R2ind29 R2ind29_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[18]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[27], x[29], x[28], x[26], x[25], x[24], x[23], x[22], x[21], x[35], x[34]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[27], x[29], x[28], x[26], x[25], x[24], x[23], x[22], x[21], x[33], x[32]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[28], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[31], x[30]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[44], x[46], x[45], x[43], x[42], x[41], x[40], x[39], x[38], x[52], x[51]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[44], x[46], x[45], x[43], x[42], x[41], x[40], x[39], x[38], x[50], x[49]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[45], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[48], x[47]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[61], x[63], x[62], x[60], x[59], x[58], x[57], x[56], x[55], x[69], x[68]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[61], x[63], x[62], x[60], x[59], x[58], x[57], x[56], x[55], x[67], x[66]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[62], x[63], x[61], x[59], x[58], x[57], x[56], x[55], x[65], x[64]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[78], x[80], x[79], x[77], x[76], x[75], x[74], x[73], x[72], x[86], x[85]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[78], x[80], x[79], x[77], x[76], x[75], x[74], x[73], x[72], x[84], x[83]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[79], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[82], x[81]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[95], x[97], x[96], x[94], x[93], x[92], x[91], x[90], x[89], x[103], x[102]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[95], x[97], x[96], x[94], x[93], x[92], x[91], x[90], x[89], x[101], x[100]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[96], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[99], x[98]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[112], x[114], x[113], x[111], x[110], x[109], x[108], x[107], x[106], x[120], x[119]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[112], x[114], x[113], x[111], x[110], x[109], x[108], x[107], x[106], x[118], x[117]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[113], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[116], x[115]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[129], x[131], x[130], x[128], x[127], x[126], x[125], x[124], x[123], x[137], x[136]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[129], x[131], x[130], x[128], x[127], x[126], x[125], x[124], x[123], x[135], x[134]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[130], x[131], x[129], x[127], x[126], x[125], x[124], x[123], x[133], x[132]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[146], x[148], x[147], x[145], x[144], x[143], x[142], x[141], x[140], x[154], x[153]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[146], x[148], x[147], x[145], x[144], x[143], x[142], x[141], x[140], x[152], x[151]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[147], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[150], x[149]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[163], x[165], x[164], x[162], x[161], x[160], x[159], x[158], x[157], x[171], x[170]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[163], x[165], x[164], x[162], x[161], x[160], x[159], x[158], x[157], x[169], x[168]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[164], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[167], x[166]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[180], x[182], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[188], x[187]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[180], x[182], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[186], x[185]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[181], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[184], x[183]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[197], x[199], x[198], x[196], x[195], x[194], x[193], x[192], x[191], x[205], x[204]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[197], x[199], x[198], x[196], x[195], x[194], x[193], x[192], x[191], x[203], x[202]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[198], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[201], x[200]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[214], x[216], x[215], x[213], x[212], x[211], x[210], x[209], x[208], x[222], x[221]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[214], x[216], x[215], x[213], x[212], x[211], x[210], x[209], x[208], x[220], x[219]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[215], x[216], x[214], x[212], x[211], x[210], x[209], x[208], x[218], x[217]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[231], x[233], x[232], x[230], x[229], x[228], x[227], x[226], x[225], x[239], x[238]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[231], x[233], x[232], x[230], x[229], x[228], x[227], x[226], x[225], x[237], x[236]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[232], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[235], x[234]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[233], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[248], x[250], x[249], x[247], x[246], x[245], x[244], x[243], x[242], x[256], x[255]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[248], x[250], x[249], x[247], x[246], x[245], x[244], x[243], x[242], x[254], x[253]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[249], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[252], x[251]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[265], x[267], x[266], x[264], x[263], x[262], x[261], x[260], x[259], x[273], x[272]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[265], x[267], x[266], x[264], x[263], x[262], x[261], x[260], x[259], x[271], x[270]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[266], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[269], x[268]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[282], x[284], x[283], x[281], x[280], x[279], x[278], x[277], x[276], x[290], x[289]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[282], x[284], x[283], x[281], x[280], x[279], x[278], x[277], x[276], x[288], x[287]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[283], x[284], x[282], x[280], x[279], x[278], x[277], x[276], x[286], x[285]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[68], x[69], x[85], x[86], x[273], x[272], x[290], x[289], x[52], x[51], x[256], x[255], x[35], x[34], x[295], x[28], x[66], x[67], x[83], x[84], x[271], x[270], x[288], x[287], x[49], x[50], x[254], x[253], x[33], x[32], x[294], x[27], x[81], x[82], x[65], x[64], x[286], x[285], x[269], x[268], x[47], x[48], x[252], x[251], x[31], x[30], x[293], x[26], x[80], x[267], x[63], x[79], x[78], x[165], x[46], x[266], x[265], x[114], x[284], x[54], x[53], x[62], x[61], x[70], x[71], x[77], x[76], x[75], x[74], x[73], x[72], x[164], x[163], x[45], x[44], x[250], x[258], x[257], x[264], x[263], x[262], x[261], x[260], x[259], x[113], x[112], x[275], x[274], x[283], x[282], x[199], x[60], x[59], x[58], x[57], x[56], x[55], x[162], x[161], x[160], x[159], x[158], x[157], x[36], x[37], x[43], x[42], x[41], x[40], x[39], x[38], x[249], x[248], x[111], x[110], x[109], x[108], x[107], x[106], x[281], x[280], x[279], x[278], x[277], x[276], x[241], x[240], x[198], x[197], x[247], x[246], x[245], x[244], x[243], x[242], x[196], x[195], x[194], x[193], x[192], x[191], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[20], x[19], x[292], x[291], x[18], x[29], x[25], x[24], x[23], x[22], x[21]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[78], x[265], x[61], x[80], x[79], x[163], x[44], x[267], x[266], x[112], x[282], x[63], x[62], x[77], x[76], x[75], x[74], x[73], x[72], x[165], x[164], x[46], x[45], x[248], x[264], x[263], x[262], x[261], x[260], x[259], x[114], x[113], x[284], x[283], x[197], x[68], x[69], x[60], x[59], x[58], x[57], x[56], x[55], x[85], x[86], x[162], x[161], x[160], x[159], x[158], x[157], x[43], x[42], x[41], x[40], x[39], x[38], x[250], x[249], x[273], x[272], x[111], x[110], x[109], x[108], x[107], x[106], x[290], x[289], x[281], x[280], x[279], x[278], x[277], x[276], x[199], x[198], x[52], x[51], x[247], x[246], x[245], x[244], x[243], x[242], x[256], x[255], x[196], x[195], x[194], x[193], x[192], x[191], x[35], x[34], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[295], x[291], x[18], x[28], x[25], x[24], x[23], x[22], x[21]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[78], x[265], x[61], x[80], x[79], x[163], x[44], x[267], x[266], x[112], x[282], x[63], x[62], x[77], x[76], x[75], x[74], x[73], x[72], x[165], x[164], x[46], x[45], x[248], x[264], x[263], x[262], x[261], x[260], x[259], x[114], x[113], x[284], x[283], x[197], x[66], x[67], x[60], x[59], x[58], x[57], x[56], x[55], x[83], x[84], x[162], x[161], x[160], x[159], x[158], x[157], x[43], x[42], x[41], x[40], x[39], x[38], x[250], x[249], x[271], x[270], x[111], x[110], x[109], x[108], x[107], x[106], x[288], x[287], x[281], x[280], x[279], x[278], x[277], x[276], x[199], x[198], x[49], x[50], x[247], x[246], x[245], x[244], x[243], x[242], x[254], x[253], x[196], x[195], x[194], x[193], x[192], x[191], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[33], x[32], x[294], x[291], x[18], x[27], x[25], x[24], x[23], x[22], x[21]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[79], x[266], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[164], x[62], x[45], x[283], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[113], x[81], x[82], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[65], x[64], x[63], x[61], x[59], x[58], x[57], x[56], x[55], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[249], x[286], x[285], x[284], x[282], x[280], x[279], x[278], x[277], x[276], x[269], x[268], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[198], x[47], x[48], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[252], x[251], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[31], x[30], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[293], x[291], x[18], x[26], x[25], x[24], x[23], x[22], x[21]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[80], x[267], x[63], x[79], x[78], x[165], x[46], x[266], x[265], x[114], x[284], x[54], x[53], x[62], x[61], x[70], x[71], x[77], x[76], x[75], x[74], x[73], x[72], x[164], x[163], x[45], x[44], x[250], x[258], x[257], x[264], x[263], x[262], x[261], x[260], x[259], x[113], x[112], x[275], x[274], x[283], x[282], x[199], x[60], x[59], x[58], x[57], x[56], x[55], x[162], x[161], x[160], x[159], x[158], x[157], x[36], x[37], x[43], x[42], x[41], x[40], x[39], x[38], x[249], x[248], x[111], x[110], x[109], x[108], x[107], x[106], x[281], x[280], x[279], x[278], x[277], x[276], x[241], x[240], x[198], x[197], x[247], x[246], x[245], x[244], x[243], x[242], x[196], x[195], x[194], x[193], x[192], x[191], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[20], x[19], x[292], x[291], x[18], x[29], x[25], x[24], x[23], x[22], x[21]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[68], x[69], x[85], x[86], x[188], x[187], x[170], x[171], x[34], x[35], x[205], x[204], x[52], x[51], x[299], x[45], x[66], x[67], x[83], x[84], x[186], x[185], x[168], x[169], x[32], x[33], x[203], x[202], x[50], x[49], x[298], x[44], x[81], x[82], x[65], x[64], x[184], x[183], x[166], x[167], x[30], x[31], x[201], x[200], x[48], x[47], x[297], x[43], x[80], x[182], x[63], x[79], x[78], x[165], x[29], x[267], x[181], x[180], x[97], x[199], x[54], x[53], x[62], x[61], x[70], x[71], x[77], x[76], x[75], x[74], x[73], x[72], x[164], x[163], x[28], x[27], x[148], x[155], x[156], x[266], x[265], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[198], x[197], x[216], x[60], x[59], x[58], x[57], x[56], x[55], x[162], x[161], x[160], x[159], x[158], x[157], x[19], x[20], x[26], x[25], x[24], x[23], x[22], x[21], x[147], x[146], x[264], x[263], x[262], x[261], x[260], x[259], x[94], x[93], x[92], x[91], x[90], x[89], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[145], x[144], x[143], x[142], x[141], x[140], x[213], x[212], x[211], x[210], x[209], x[208], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[37], x[36], x[296], x[291], x[18], x[46], x[42], x[41], x[40], x[39], x[38]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[78], x[180], x[61], x[80], x[79], x[163], x[27], x[182], x[181], x[95], x[265], x[197], x[63], x[62], x[77], x[76], x[75], x[74], x[73], x[72], x[165], x[164], x[29], x[28], x[146], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[267], x[266], x[199], x[198], x[214], x[68], x[69], x[60], x[59], x[58], x[57], x[56], x[55], x[85], x[86], x[162], x[161], x[160], x[159], x[158], x[157], x[26], x[25], x[24], x[23], x[22], x[21], x[148], x[147], x[188], x[187], x[94], x[93], x[92], x[91], x[90], x[89], x[170], x[171], x[264], x[263], x[262], x[261], x[260], x[259], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[34], x[35], x[145], x[144], x[143], x[142], x[141], x[140], x[205], x[204], x[213], x[212], x[211], x[210], x[209], x[208], x[52], x[51], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[299], x[291], x[18], x[45], x[42], x[41], x[40], x[39], x[38]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[78], x[180], x[61], x[80], x[79], x[163], x[27], x[182], x[181], x[95], x[265], x[197], x[63], x[62], x[77], x[76], x[75], x[74], x[73], x[72], x[165], x[164], x[29], x[28], x[146], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[267], x[266], x[199], x[198], x[214], x[66], x[67], x[60], x[59], x[58], x[57], x[56], x[55], x[83], x[84], x[162], x[161], x[160], x[159], x[158], x[157], x[26], x[25], x[24], x[23], x[22], x[21], x[148], x[147], x[186], x[185], x[94], x[93], x[92], x[91], x[90], x[89], x[168], x[169], x[264], x[263], x[262], x[261], x[260], x[259], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[32], x[33], x[145], x[144], x[143], x[142], x[141], x[140], x[203], x[202], x[213], x[212], x[211], x[210], x[209], x[208], x[50], x[49], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[298], x[291], x[18], x[44], x[42], x[41], x[40], x[39], x[38]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[79], x[181], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[164], x[62], x[28], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[96], x[266], x[198], x[81], x[82], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[65], x[64], x[63], x[61], x[59], x[58], x[57], x[56], x[55], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[147], x[184], x[183], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[166], x[167], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[215], x[30], x[31], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[201], x[200], x[216], x[214], x[212], x[211], x[210], x[209], x[208], x[48], x[47], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[297], x[291], x[18], x[43], x[42], x[41], x[40], x[39], x[38]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[80], x[182], x[63], x[79], x[78], x[165], x[29], x[267], x[181], x[180], x[97], x[199], x[54], x[53], x[62], x[61], x[70], x[71], x[77], x[76], x[75], x[74], x[73], x[72], x[164], x[163], x[28], x[27], x[148], x[155], x[156], x[266], x[265], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[198], x[197], x[216], x[60], x[59], x[58], x[57], x[56], x[55], x[162], x[161], x[160], x[159], x[158], x[157], x[19], x[20], x[26], x[25], x[24], x[23], x[22], x[21], x[147], x[146], x[264], x[263], x[262], x[261], x[260], x[259], x[94], x[93], x[92], x[91], x[90], x[89], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[145], x[144], x[143], x[142], x[141], x[140], x[213], x[212], x[211], x[210], x[209], x[208], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[37], x[36], x[296], x[291], x[18], x[46], x[42], x[41], x[40], x[39], x[38]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[52], x[51], x[34], x[35], x[85], x[86], x[69], x[68], x[303], x[62], x[49], x[50], x[32], x[33], x[83], x[84], x[67], x[66], x[302], x[61], x[47], x[48], x[30], x[31], x[81], x[82], x[65], x[64], x[301], x[60], x[29], x[46], x[28], x[27], x[148], x[45], x[44], x[250], x[80], x[19], x[20], x[26], x[25], x[24], x[23], x[22], x[21], x[147], x[146], x[36], x[37], x[43], x[42], x[41], x[40], x[39], x[38], x[249], x[248], x[79], x[78], x[165], x[145], x[144], x[143], x[142], x[141], x[140], x[247], x[246], x[245], x[244], x[243], x[242], x[70], x[71], x[77], x[76], x[75], x[74], x[73], x[72], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[54], x[53], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[300], x[291], x[18], x[63], x[59], x[58], x[57], x[56], x[55]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[44], x[27], x[46], x[45], x[248], x[29], x[28], x[146], x[78], x[43], x[42], x[41], x[40], x[39], x[38], x[250], x[249], x[26], x[25], x[24], x[23], x[22], x[21], x[148], x[147], x[80], x[79], x[163], x[52], x[51], x[247], x[246], x[245], x[244], x[243], x[242], x[34], x[35], x[145], x[144], x[143], x[142], x[141], x[140], x[77], x[76], x[75], x[74], x[73], x[72], x[165], x[164], x[85], x[86], x[162], x[161], x[160], x[159], x[158], x[157], x[69], x[68], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[303], x[291], x[18], x[62], x[59], x[58], x[57], x[56], x[55]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[44], x[27], x[46], x[45], x[248], x[29], x[28], x[146], x[78], x[43], x[42], x[41], x[40], x[39], x[38], x[250], x[249], x[26], x[25], x[24], x[23], x[22], x[21], x[148], x[147], x[80], x[79], x[163], x[49], x[50], x[247], x[246], x[245], x[244], x[243], x[242], x[32], x[33], x[145], x[144], x[143], x[142], x[141], x[140], x[77], x[76], x[75], x[74], x[73], x[72], x[165], x[164], x[83], x[84], x[162], x[161], x[160], x[159], x[158], x[157], x[67], x[66], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[302], x[291], x[18], x[61], x[59], x[58], x[57], x[56], x[55]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[45], x[28], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[249], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[147], x[79], x[47], x[48], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[30], x[31], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[164], x[81], x[82], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[65], x[64], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[301], x[291], x[18], x[60], x[59], x[58], x[57], x[56], x[55]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[29], x[46], x[28], x[27], x[148], x[45], x[44], x[250], x[80], x[19], x[20], x[26], x[25], x[24], x[23], x[22], x[21], x[147], x[146], x[36], x[37], x[43], x[42], x[41], x[40], x[39], x[38], x[249], x[248], x[79], x[78], x[165], x[145], x[144], x[143], x[142], x[141], x[140], x[247], x[246], x[245], x[244], x[243], x[242], x[70], x[71], x[77], x[76], x[75], x[74], x[73], x[72], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[54], x[53], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[300], x[291], x[18], x[63], x[59], x[58], x[57], x[56], x[55]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[52], x[51], x[34], x[35], x[136], x[137], x[153], x[154], x[68], x[69], x[102], x[103], x[86], x[85], x[307], x[79], x[49], x[50], x[32], x[33], x[134], x[135], x[151], x[152], x[66], x[67], x[100], x[101], x[84], x[83], x[306], x[78], x[47], x[48], x[30], x[31], x[149], x[150], x[132], x[133], x[65], x[64], x[98], x[99], x[82], x[81], x[305], x[77], x[29], x[46], x[28], x[27], x[148], x[45], x[44], x[250], x[233], x[131], x[97], x[19], x[20], x[26], x[25], x[24], x[23], x[22], x[21], x[147], x[146], x[36], x[37], x[43], x[42], x[41], x[40], x[39], x[38], x[249], x[248], x[63], x[121], x[122], x[232], x[231], x[138], x[139], x[130], x[129], x[96], x[95], x[182], x[145], x[144], x[143], x[142], x[141], x[140], x[247], x[246], x[245], x[244], x[243], x[242], x[54], x[53], x[62], x[61], x[230], x[229], x[228], x[227], x[226], x[225], x[128], x[127], x[126], x[125], x[124], x[123], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[60], x[59], x[58], x[57], x[56], x[55], x[179], x[178], x[177], x[176], x[175], x[174], x[71], x[70], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[304], x[291], x[18], x[80], x[76], x[75], x[74], x[73], x[72]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[44], x[27], x[46], x[45], x[248], x[29], x[28], x[146], x[231], x[129], x[95], x[43], x[42], x[41], x[40], x[39], x[38], x[250], x[249], x[26], x[25], x[24], x[23], x[22], x[21], x[148], x[147], x[61], x[233], x[232], x[131], x[130], x[97], x[96], x[180], x[52], x[51], x[247], x[246], x[245], x[244], x[243], x[242], x[34], x[35], x[145], x[144], x[143], x[142], x[141], x[140], x[63], x[62], x[136], x[137], x[230], x[229], x[228], x[227], x[226], x[225], x[153], x[154], x[128], x[127], x[126], x[125], x[124], x[123], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[68], x[69], x[60], x[59], x[58], x[57], x[56], x[55], x[102], x[103], x[179], x[178], x[177], x[176], x[175], x[174], x[86], x[85], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[307], x[291], x[18], x[79], x[76], x[75], x[74], x[73], x[72]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[44], x[27], x[46], x[45], x[248], x[29], x[28], x[146], x[231], x[129], x[95], x[43], x[42], x[41], x[40], x[39], x[38], x[250], x[249], x[26], x[25], x[24], x[23], x[22], x[21], x[148], x[147], x[61], x[233], x[232], x[131], x[130], x[97], x[96], x[180], x[49], x[50], x[247], x[246], x[245], x[244], x[243], x[242], x[32], x[33], x[145], x[144], x[143], x[142], x[141], x[140], x[63], x[62], x[134], x[135], x[230], x[229], x[228], x[227], x[226], x[225], x[151], x[152], x[128], x[127], x[126], x[125], x[124], x[123], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[66], x[67], x[60], x[59], x[58], x[57], x[56], x[55], x[100], x[101], x[179], x[178], x[177], x[176], x[175], x[174], x[84], x[83], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[306], x[291], x[18], x[78], x[76], x[75], x[74], x[73], x[72]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[45], x[28], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[249], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[147], x[130], x[232], x[96], x[47], x[48], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[30], x[31], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[62], x[149], x[150], x[131], x[129], x[127], x[126], x[125], x[124], x[123], x[132], x[133], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[181], x[65], x[64], x[63], x[61], x[59], x[58], x[57], x[56], x[55], x[98], x[99], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[82], x[81], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[305], x[291], x[18], x[77], x[76], x[75], x[74], x[73], x[72]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[29], x[46], x[28], x[27], x[148], x[45], x[44], x[250], x[233], x[131], x[97], x[19], x[20], x[26], x[25], x[24], x[23], x[22], x[21], x[147], x[146], x[36], x[37], x[43], x[42], x[41], x[40], x[39], x[38], x[249], x[248], x[63], x[121], x[122], x[232], x[231], x[138], x[139], x[130], x[129], x[96], x[95], x[182], x[145], x[144], x[143], x[142], x[141], x[140], x[247], x[246], x[245], x[244], x[243], x[242], x[54], x[53], x[62], x[61], x[230], x[229], x[228], x[227], x[226], x[225], x[128], x[127], x[126], x[125], x[124], x[123], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[60], x[59], x[58], x[57], x[56], x[55], x[179], x[178], x[177], x[176], x[175], x[174], x[71], x[70], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[304], x[291], x[18], x[80], x[76], x[75], x[74], x[73], x[72]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[136], x[137], x[153], x[154], x[205], x[204], x[222], x[221], x[119], x[120], x[170], x[171], x[103], x[102], x[311], x[96], x[134], x[135], x[151], x[152], x[203], x[202], x[220], x[219], x[117], x[118], x[168], x[169], x[101], x[100], x[310], x[95], x[149], x[150], x[132], x[133], x[218], x[217], x[201], x[200], x[115], x[116], x[166], x[167], x[99], x[98], x[309], x[94], x[148], x[199], x[233], x[147], x[146], x[131], x[114], x[198], x[197], x[216], x[46], x[165], x[121], x[122], x[232], x[231], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[113], x[112], x[80], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[207], x[206], x[45], x[44], x[164], x[163], x[267], x[230], x[229], x[228], x[227], x[226], x[225], x[128], x[127], x[126], x[125], x[124], x[123], x[104], x[105], x[111], x[110], x[109], x[108], x[107], x[106], x[79], x[78], x[213], x[212], x[211], x[210], x[209], x[208], x[43], x[42], x[41], x[40], x[39], x[38], x[155], x[156], x[162], x[161], x[160], x[159], x[158], x[157], x[266], x[265], x[77], x[76], x[75], x[74], x[73], x[72], x[264], x[263], x[262], x[261], x[260], x[259], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[88], x[87], x[308], x[291], x[18], x[97], x[93], x[92], x[91], x[90], x[89]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[146], x[197], x[231], x[148], x[147], x[129], x[112], x[199], x[198], x[214], x[44], x[163], x[233], x[232], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[114], x[113], x[78], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[46], x[45], x[165], x[164], x[265], x[136], x[137], x[230], x[229], x[228], x[227], x[226], x[225], x[153], x[154], x[128], x[127], x[126], x[125], x[124], x[123], x[111], x[110], x[109], x[108], x[107], x[106], x[80], x[79], x[205], x[204], x[213], x[212], x[211], x[210], x[209], x[208], x[222], x[221], x[43], x[42], x[41], x[40], x[39], x[38], x[162], x[161], x[160], x[159], x[158], x[157], x[267], x[266], x[119], x[120], x[77], x[76], x[75], x[74], x[73], x[72], x[170], x[171], x[264], x[263], x[262], x[261], x[260], x[259], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[103], x[102], x[311], x[291], x[18], x[96], x[93], x[92], x[91], x[90], x[89]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[146], x[197], x[231], x[148], x[147], x[129], x[112], x[199], x[198], x[214], x[44], x[163], x[233], x[232], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[114], x[113], x[78], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[46], x[45], x[165], x[164], x[265], x[134], x[135], x[230], x[229], x[228], x[227], x[226], x[225], x[151], x[152], x[128], x[127], x[126], x[125], x[124], x[123], x[111], x[110], x[109], x[108], x[107], x[106], x[80], x[79], x[203], x[202], x[213], x[212], x[211], x[210], x[209], x[208], x[220], x[219], x[43], x[42], x[41], x[40], x[39], x[38], x[162], x[161], x[160], x[159], x[158], x[157], x[267], x[266], x[117], x[118], x[77], x[76], x[75], x[74], x[73], x[72], x[168], x[169], x[264], x[263], x[262], x[261], x[260], x[259], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[101], x[100], x[310], x[291], x[18], x[95], x[93], x[92], x[91], x[90], x[89]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[147], x[198], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[130], x[232], x[113], x[45], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[215], x[164], x[149], x[150], x[131], x[129], x[127], x[126], x[125], x[124], x[123], x[132], x[133], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[79], x[218], x[217], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[201], x[200], x[216], x[214], x[212], x[211], x[210], x[209], x[208], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[266], x[115], x[116], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[166], x[167], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[99], x[98], x[309], x[291], x[18], x[94], x[93], x[92], x[91], x[90], x[89]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[148], x[199], x[233], x[147], x[146], x[131], x[114], x[198], x[197], x[216], x[46], x[165], x[121], x[122], x[232], x[231], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[113], x[112], x[80], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[207], x[206], x[45], x[44], x[164], x[163], x[267], x[230], x[229], x[228], x[227], x[226], x[225], x[128], x[127], x[126], x[125], x[124], x[123], x[104], x[105], x[111], x[110], x[109], x[108], x[107], x[106], x[79], x[78], x[213], x[212], x[211], x[210], x[209], x[208], x[43], x[42], x[41], x[40], x[39], x[38], x[155], x[156], x[162], x[161], x[160], x[159], x[158], x[157], x[266], x[265], x[77], x[76], x[75], x[74], x[73], x[72], x[264], x[263], x[262], x[261], x[260], x[259], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[88], x[87], x[308], x[291], x[18], x[97], x[93], x[92], x[91], x[90], x[89]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[136], x[137], x[153], x[154], x[256], x[255], x[239], x[238], x[102], x[103], x[290], x[289], x[120], x[119], x[315], x[113], x[134], x[135], x[151], x[152], x[254], x[253], x[237], x[236], x[100], x[101], x[288], x[287], x[118], x[117], x[314], x[112], x[149], x[150], x[132], x[133], x[252], x[251], x[235], x[234], x[98], x[99], x[286], x[285], x[116], x[115], x[313], x[111], x[148], x[250], x[233], x[147], x[146], x[131], x[97], x[29], x[249], x[248], x[199], x[121], x[122], x[232], x[231], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[96], x[95], x[182], x[224], x[223], x[28], x[27], x[241], x[240], x[247], x[246], x[245], x[244], x[243], x[242], x[198], x[197], x[284], x[230], x[229], x[228], x[227], x[226], x[225], x[128], x[127], x[126], x[125], x[124], x[123], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[26], x[25], x[24], x[23], x[22], x[21], x[196], x[195], x[194], x[193], x[192], x[191], x[275], x[274], x[283], x[282], x[179], x[178], x[177], x[176], x[175], x[174], x[281], x[280], x[279], x[278], x[277], x[276], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[105], x[104], x[312], x[291], x[18], x[114], x[110], x[109], x[108], x[107], x[106]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[146], x[248], x[231], x[148], x[147], x[129], x[95], x[250], x[249], x[197], x[27], x[233], x[232], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[97], x[96], x[180], x[247], x[246], x[245], x[244], x[243], x[242], x[199], x[198], x[29], x[28], x[282], x[136], x[137], x[230], x[229], x[228], x[227], x[226], x[225], x[153], x[154], x[128], x[127], x[126], x[125], x[124], x[123], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[256], x[255], x[196], x[195], x[194], x[193], x[192], x[191], x[239], x[238], x[26], x[25], x[24], x[23], x[22], x[21], x[284], x[283], x[102], x[103], x[179], x[178], x[177], x[176], x[175], x[174], x[290], x[289], x[281], x[280], x[279], x[278], x[277], x[276], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[120], x[119], x[315], x[291], x[18], x[113], x[110], x[109], x[108], x[107], x[106]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[146], x[248], x[231], x[148], x[147], x[129], x[95], x[250], x[249], x[197], x[27], x[233], x[232], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[97], x[96], x[180], x[247], x[246], x[245], x[244], x[243], x[242], x[199], x[198], x[29], x[28], x[282], x[134], x[135], x[230], x[229], x[228], x[227], x[226], x[225], x[151], x[152], x[128], x[127], x[126], x[125], x[124], x[123], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[254], x[253], x[196], x[195], x[194], x[193], x[192], x[191], x[237], x[236], x[26], x[25], x[24], x[23], x[22], x[21], x[284], x[283], x[100], x[101], x[179], x[178], x[177], x[176], x[175], x[174], x[288], x[287], x[281], x[280], x[279], x[278], x[277], x[276], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[118], x[117], x[314], x[291], x[18], x[112], x[110], x[109], x[108], x[107], x[106]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[147], x[249], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[130], x[232], x[96], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[198], x[28], x[149], x[150], x[131], x[129], x[127], x[126], x[125], x[124], x[123], x[132], x[133], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[181], x[252], x[251], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[235], x[234], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[283], x[98], x[99], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[286], x[285], x[284], x[282], x[280], x[279], x[278], x[277], x[276], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[116], x[115], x[313], x[291], x[18], x[111], x[110], x[109], x[108], x[107], x[106]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[148], x[250], x[233], x[147], x[146], x[131], x[97], x[29], x[249], x[248], x[199], x[121], x[122], x[232], x[231], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[96], x[95], x[182], x[224], x[223], x[28], x[27], x[241], x[240], x[247], x[246], x[245], x[244], x[243], x[242], x[198], x[197], x[284], x[230], x[229], x[228], x[227], x[226], x[225], x[128], x[127], x[126], x[125], x[124], x[123], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[26], x[25], x[24], x[23], x[22], x[21], x[196], x[195], x[194], x[193], x[192], x[191], x[275], x[274], x[283], x[282], x[179], x[178], x[177], x[176], x[175], x[174], x[281], x[280], x[279], x[278], x[277], x[276], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[105], x[104], x[312], x[291], x[18], x[114], x[110], x[109], x[108], x[107], x[106]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[119], x[120], x[102], x[103], x[153], x[154], x[137], x[136], x[319], x[117], x[118], x[100], x[101], x[151], x[152], x[135], x[134], x[318], x[115], x[116], x[98], x[99], x[149], x[150], x[133], x[132], x[317], x[97], x[114], x[148], x[96], x[95], x[182], x[113], x[112], x[80], x[147], x[146], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[104], x[105], x[111], x[110], x[109], x[108], x[107], x[106], x[79], x[78], x[233], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[179], x[178], x[177], x[176], x[175], x[174], x[77], x[76], x[75], x[74], x[73], x[72], x[232], x[231], x[128], x[230], x[229], x[228], x[227], x[226], x[225], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[122], x[121], x[316], x[291], x[18], x[131], x[127], x[126], x[125], x[124], x[123]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[112], x[95], x[146], x[114], x[113], x[78], x[97], x[96], x[180], x[148], x[147], x[129], x[111], x[110], x[109], x[108], x[107], x[106], x[80], x[79], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[231], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[119], x[120], x[77], x[76], x[75], x[74], x[73], x[72], x[102], x[103], x[179], x[178], x[177], x[176], x[175], x[174], x[233], x[232], x[153], x[154], x[128], x[230], x[229], x[228], x[227], x[226], x[225], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[137], x[136], x[319], x[291], x[18], x[130], x[127], x[126], x[125], x[124], x[123]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[112], x[95], x[146], x[114], x[113], x[78], x[97], x[96], x[180], x[148], x[147], x[111], x[110], x[109], x[108], x[107], x[106], x[80], x[79], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[231], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[117], x[118], x[77], x[76], x[75], x[74], x[73], x[72], x[100], x[101], x[179], x[178], x[177], x[176], x[175], x[174], x[233], x[232], x[151], x[152], x[128], x[230], x[229], x[228], x[227], x[226], x[225], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[135], x[134], x[318], x[291], x[18], x[129], x[127], x[126], x[125], x[124], x[123]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[113], x[96], x[147], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[79], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[181], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[130], x[115], x[116], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[98], x[99], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[232], x[149], x[150], x[131], x[129], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[133], x[132], x[317], x[291], x[18], x[128], x[127], x[126], x[125], x[124], x[123]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[97], x[114], x[148], x[96], x[95], x[182], x[113], x[112], x[80], x[147], x[146], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[104], x[105], x[111], x[110], x[109], x[108], x[107], x[106], x[79], x[78], x[233], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[179], x[178], x[177], x[176], x[175], x[174], x[77], x[76], x[75], x[74], x[73], x[72], x[232], x[231], x[128], x[230], x[229], x[228], x[227], x[226], x[225], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[122], x[121], x[316], x[291], x[18], x[131], x[127], x[126], x[125], x[124], x[123]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[119], x[120], x[102], x[103], x[68], x[69], x[85], x[86], x[136], x[137], x[52], x[51], x[154], x[153], x[323], x[147], x[117], x[118], x[100], x[101], x[66], x[67], x[83], x[84], x[134], x[135], x[49], x[50], x[152], x[151], x[322], x[146], x[115], x[116], x[98], x[99], x[81], x[82], x[65], x[64], x[132], x[133], x[47], x[48], x[150], x[149], x[321], x[145], x[97], x[114], x[96], x[95], x[182], x[113], x[112], x[80], x[131], x[63], x[165], x[46], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[104], x[105], x[111], x[110], x[109], x[108], x[107], x[106], x[79], x[78], x[130], x[129], x[233], x[54], x[53], x[62], x[61], x[70], x[71], x[164], x[163], x[45], x[44], x[250], x[179], x[178], x[177], x[176], x[175], x[174], x[77], x[76], x[75], x[74], x[73], x[72], x[121], x[122], x[128], x[127], x[126], x[125], x[124], x[123], x[232], x[231], x[60], x[59], x[58], x[57], x[56], x[55], x[162], x[161], x[160], x[159], x[158], x[157], x[36], x[37], x[43], x[42], x[41], x[40], x[39], x[38], x[249], x[248], x[230], x[229], x[228], x[227], x[226], x[225], x[247], x[246], x[245], x[244], x[243], x[242], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[139], x[138], x[320], x[291], x[18], x[148], x[144], x[143], x[142], x[141], x[140]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[112], x[95], x[114], x[113], x[78], x[97], x[96], x[180], x[129], x[61], x[163], x[44], x[111], x[110], x[109], x[108], x[107], x[106], x[80], x[79], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[131], x[130], x[231], x[63], x[62], x[165], x[164], x[46], x[45], x[248], x[119], x[120], x[77], x[76], x[75], x[74], x[73], x[72], x[102], x[103], x[179], x[178], x[177], x[176], x[175], x[174], x[128], x[127], x[126], x[125], x[124], x[123], x[233], x[232], x[68], x[69], x[60], x[59], x[58], x[57], x[56], x[55], x[85], x[86], x[162], x[161], x[160], x[159], x[158], x[157], x[43], x[42], x[41], x[40], x[39], x[38], x[250], x[249], x[136], x[137], x[230], x[229], x[228], x[227], x[226], x[225], x[52], x[51], x[247], x[246], x[245], x[244], x[243], x[242], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[154], x[153], x[323], x[291], x[18], x[147], x[144], x[143], x[142], x[141], x[140]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[112], x[95], x[114], x[113], x[78], x[97], x[96], x[180], x[129], x[61], x[163], x[44], x[111], x[110], x[109], x[108], x[107], x[106], x[80], x[79], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[131], x[130], x[231], x[63], x[62], x[165], x[164], x[46], x[45], x[248], x[117], x[118], x[77], x[76], x[75], x[74], x[73], x[72], x[100], x[101], x[179], x[178], x[177], x[176], x[175], x[174], x[128], x[127], x[126], x[125], x[124], x[123], x[233], x[232], x[66], x[67], x[60], x[59], x[58], x[57], x[56], x[55], x[83], x[84], x[162], x[161], x[160], x[159], x[158], x[157], x[43], x[42], x[41], x[40], x[39], x[38], x[250], x[249], x[134], x[135], x[230], x[229], x[228], x[227], x[226], x[225], x[49], x[50], x[247], x[246], x[245], x[244], x[243], x[242], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[152], x[151], x[322], x[291], x[18], x[146], x[144], x[143], x[142], x[141], x[140]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[113], x[96], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[79], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[181], x[130], x[164], x[62], x[45], x[115], x[116], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[98], x[99], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[131], x[129], x[127], x[126], x[125], x[124], x[123], x[232], x[81], x[82], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[65], x[64], x[63], x[61], x[59], x[58], x[57], x[56], x[55], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[249], x[132], x[133], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[47], x[48], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[150], x[149], x[321], x[291], x[18], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[97], x[114], x[96], x[95], x[182], x[113], x[112], x[80], x[131], x[63], x[165], x[46], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[104], x[105], x[111], x[110], x[109], x[108], x[107], x[106], x[79], x[78], x[130], x[129], x[233], x[54], x[53], x[62], x[61], x[70], x[71], x[164], x[163], x[45], x[44], x[250], x[179], x[178], x[177], x[176], x[175], x[174], x[77], x[76], x[75], x[74], x[73], x[72], x[121], x[122], x[128], x[127], x[126], x[125], x[124], x[123], x[232], x[231], x[60], x[59], x[58], x[57], x[56], x[55], x[162], x[161], x[160], x[159], x[158], x[157], x[36], x[37], x[43], x[42], x[41], x[40], x[39], x[38], x[249], x[248], x[230], x[229], x[228], x[227], x[226], x[225], x[247], x[246], x[245], x[244], x[243], x[242], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[139], x[138], x[320], x[291], x[18], x[148], x[144], x[143], x[142], x[141], x[140]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[205], x[204], x[222], x[221], x[52], x[51], x[34], x[35], x[188], x[187], x[68], x[69], x[171], x[170], x[327], x[164], x[203], x[202], x[220], x[219], x[49], x[50], x[32], x[33], x[186], x[185], x[66], x[67], x[169], x[168], x[326], x[163], x[218], x[217], x[201], x[200], x[47], x[48], x[30], x[31], x[184], x[183], x[65], x[64], x[167], x[166], x[325], x[162], x[199], x[29], x[198], x[197], x[216], x[46], x[182], x[28], x[27], x[148], x[250], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[207], x[206], x[45], x[44], x[181], x[180], x[97], x[19], x[20], x[26], x[25], x[24], x[23], x[22], x[21], x[147], x[146], x[36], x[37], x[249], x[248], x[63], x[213], x[212], x[211], x[210], x[209], x[208], x[43], x[42], x[41], x[40], x[39], x[38], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[145], x[144], x[143], x[142], x[141], x[140], x[247], x[246], x[245], x[244], x[243], x[242], x[54], x[53], x[62], x[61], x[94], x[93], x[92], x[91], x[90], x[89], x[60], x[59], x[58], x[57], x[56], x[55], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[156], x[155], x[324], x[291], x[18], x[165], x[161], x[160], x[159], x[158], x[157]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[197], x[27], x[199], x[198], x[214], x[44], x[180], x[248], x[29], x[28], x[146], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[46], x[45], x[182], x[181], x[95], x[250], x[249], x[26], x[25], x[24], x[23], x[22], x[21], x[148], x[147], x[61], x[205], x[204], x[213], x[212], x[211], x[210], x[209], x[208], x[222], x[221], x[43], x[42], x[41], x[40], x[39], x[38], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[52], x[51], x[247], x[246], x[245], x[244], x[243], x[242], x[34], x[35], x[145], x[144], x[143], x[142], x[141], x[140], x[63], x[62], x[188], x[187], x[94], x[93], x[92], x[91], x[90], x[89], x[68], x[69], x[60], x[59], x[58], x[57], x[56], x[55], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[171], x[170], x[327], x[291], x[18], x[164], x[161], x[160], x[159], x[158], x[157]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[197], x[27], x[199], x[198], x[214], x[44], x[180], x[248], x[29], x[28], x[146], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[46], x[45], x[182], x[181], x[95], x[250], x[249], x[26], x[25], x[24], x[23], x[22], x[21], x[148], x[147], x[61], x[203], x[202], x[213], x[212], x[211], x[210], x[209], x[208], x[220], x[219], x[43], x[42], x[41], x[40], x[39], x[38], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[49], x[50], x[247], x[246], x[245], x[244], x[243], x[242], x[32], x[33], x[145], x[144], x[143], x[142], x[141], x[140], x[63], x[62], x[186], x[185], x[94], x[93], x[92], x[91], x[90], x[89], x[66], x[67], x[60], x[59], x[58], x[57], x[56], x[55], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[169], x[168], x[326], x[291], x[18], x[163], x[161], x[160], x[159], x[158], x[157]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[198], x[28], x[45], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[215], x[181], x[249], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[147], x[218], x[217], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[201], x[200], x[216], x[214], x[212], x[211], x[210], x[209], x[208], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[96], x[47], x[48], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[30], x[31], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[62], x[184], x[183], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[65], x[64], x[63], x[61], x[59], x[58], x[57], x[56], x[55], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[167], x[166], x[325], x[291], x[18], x[162], x[161], x[160], x[159], x[158], x[157]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[199], x[29], x[198], x[197], x[216], x[46], x[182], x[28], x[27], x[148], x[250], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[207], x[206], x[45], x[44], x[181], x[180], x[97], x[19], x[20], x[26], x[25], x[24], x[23], x[22], x[21], x[147], x[146], x[36], x[37], x[249], x[248], x[63], x[213], x[212], x[211], x[210], x[209], x[208], x[43], x[42], x[41], x[40], x[39], x[38], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[145], x[144], x[143], x[142], x[141], x[140], x[247], x[246], x[245], x[244], x[243], x[242], x[54], x[53], x[62], x[61], x[94], x[93], x[92], x[91], x[90], x[89], x[60], x[59], x[58], x[57], x[56], x[55], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[156], x[155], x[324], x[291], x[18], x[165], x[161], x[160], x[159], x[158], x[157]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[205], x[204], x[222], x[221], x[136], x[137], x[153], x[154], x[170], x[171], x[119], x[120], x[188], x[187], x[331], x[181], x[203], x[202], x[220], x[219], x[134], x[135], x[151], x[152], x[168], x[169], x[117], x[118], x[186], x[185], x[330], x[180], x[218], x[217], x[201], x[200], x[149], x[150], x[132], x[133], x[166], x[167], x[115], x[116], x[184], x[183], x[329], x[179], x[199], x[148], x[198], x[197], x[216], x[46], x[165], x[233], x[147], x[146], x[131], x[114], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[207], x[206], x[45], x[44], x[164], x[163], x[267], x[121], x[122], x[232], x[231], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[113], x[112], x[80], x[213], x[212], x[211], x[210], x[209], x[208], x[43], x[42], x[41], x[40], x[39], x[38], x[155], x[156], x[162], x[161], x[160], x[159], x[158], x[157], x[266], x[265], x[230], x[229], x[228], x[227], x[226], x[225], x[128], x[127], x[126], x[125], x[124], x[123], x[104], x[105], x[111], x[110], x[109], x[108], x[107], x[106], x[79], x[78], x[264], x[263], x[262], x[261], x[260], x[259], x[77], x[76], x[75], x[74], x[73], x[72], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[173], x[172], x[328], x[291], x[18], x[182], x[178], x[177], x[176], x[175], x[174]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[197], x[146], x[199], x[198], x[214], x[44], x[163], x[231], x[148], x[147], x[129], x[112], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[46], x[45], x[165], x[164], x[265], x[233], x[232], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[114], x[113], x[78], x[205], x[204], x[213], x[212], x[211], x[210], x[209], x[208], x[222], x[221], x[43], x[42], x[41], x[40], x[39], x[38], x[162], x[161], x[160], x[159], x[158], x[157], x[267], x[266], x[136], x[137], x[230], x[229], x[228], x[227], x[226], x[225], x[153], x[154], x[128], x[127], x[126], x[125], x[124], x[123], x[111], x[110], x[109], x[108], x[107], x[106], x[80], x[79], x[170], x[171], x[264], x[263], x[262], x[261], x[260], x[259], x[119], x[120], x[77], x[76], x[75], x[74], x[73], x[72], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[188], x[187], x[331], x[291], x[18], x[181], x[178], x[177], x[176], x[175], x[174]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[197], x[146], x[199], x[198], x[214], x[44], x[163], x[231], x[148], x[147], x[129], x[112], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[46], x[45], x[165], x[164], x[265], x[233], x[232], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[114], x[113], x[78], x[203], x[202], x[213], x[212], x[211], x[210], x[209], x[208], x[220], x[219], x[43], x[42], x[41], x[40], x[39], x[38], x[162], x[161], x[160], x[159], x[158], x[157], x[267], x[266], x[134], x[135], x[230], x[229], x[228], x[227], x[226], x[225], x[151], x[152], x[128], x[127], x[126], x[125], x[124], x[123], x[111], x[110], x[109], x[108], x[107], x[106], x[80], x[79], x[168], x[169], x[264], x[263], x[262], x[261], x[260], x[259], x[117], x[118], x[77], x[76], x[75], x[74], x[73], x[72], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[186], x[185], x[330], x[291], x[18], x[180], x[178], x[177], x[176], x[175], x[174]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[198], x[147], x[45], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[215], x[164], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[130], x[232], x[113], x[218], x[217], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[201], x[200], x[216], x[214], x[212], x[211], x[210], x[209], x[208], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[266], x[149], x[150], x[131], x[129], x[127], x[126], x[125], x[124], x[123], x[132], x[133], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[79], x[166], x[167], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[115], x[116], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[184], x[183], x[329], x[291], x[18], x[179], x[178], x[177], x[176], x[175], x[174]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[199], x[148], x[198], x[197], x[216], x[46], x[165], x[233], x[147], x[146], x[131], x[114], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[207], x[206], x[45], x[44], x[164], x[163], x[267], x[121], x[122], x[232], x[231], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[113], x[112], x[80], x[213], x[212], x[211], x[210], x[209], x[208], x[43], x[42], x[41], x[40], x[39], x[38], x[155], x[156], x[162], x[161], x[160], x[159], x[158], x[157], x[266], x[265], x[230], x[229], x[228], x[227], x[226], x[225], x[128], x[127], x[126], x[125], x[124], x[123], x[104], x[105], x[111], x[110], x[109], x[108], x[107], x[106], x[79], x[78], x[264], x[263], x[262], x[261], x[260], x[259], x[77], x[76], x[75], x[74], x[73], x[72], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[173], x[172], x[328], x[291], x[18], x[182], x[178], x[177], x[176], x[175], x[174]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[188], x[187], x[170], x[171], x[273], x[272], x[290], x[289], x[222], x[221], x[239], x[238], x[205], x[204], x[335], x[198], x[186], x[185], x[168], x[169], x[271], x[270], x[288], x[287], x[220], x[219], x[237], x[236], x[203], x[202], x[334], x[197], x[184], x[183], x[166], x[167], x[286], x[285], x[269], x[268], x[218], x[217], x[235], x[234], x[201], x[200], x[333], x[196], x[165], x[182], x[164], x[163], x[267], x[181], x[180], x[97], x[216], x[114], x[284], x[233], x[155], x[156], x[162], x[161], x[160], x[159], x[158], x[157], x[266], x[265], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[215], x[214], x[46], x[258], x[257], x[113], x[112], x[275], x[274], x[283], x[282], x[232], x[231], x[29], x[264], x[263], x[262], x[261], x[260], x[259], x[94], x[93], x[92], x[91], x[90], x[89], x[207], x[206], x[213], x[212], x[211], x[210], x[209], x[208], x[45], x[44], x[111], x[110], x[109], x[108], x[107], x[106], x[281], x[280], x[279], x[278], x[277], x[276], x[224], x[223], x[230], x[229], x[228], x[227], x[226], x[225], x[28], x[27], x[43], x[42], x[41], x[40], x[39], x[38], x[26], x[25], x[24], x[23], x[22], x[21], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[190], x[189], x[332], x[291], x[18], x[199], x[195], x[194], x[193], x[192], x[191]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[180], x[163], x[182], x[181], x[95], x[165], x[164], x[265], x[214], x[112], x[282], x[231], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[162], x[161], x[160], x[159], x[158], x[157], x[267], x[266], x[216], x[215], x[44], x[114], x[113], x[284], x[283], x[233], x[232], x[27], x[188], x[187], x[94], x[93], x[92], x[91], x[90], x[89], x[170], x[171], x[264], x[263], x[262], x[261], x[260], x[259], x[213], x[212], x[211], x[210], x[209], x[208], x[46], x[45], x[273], x[272], x[111], x[110], x[109], x[108], x[107], x[106], x[290], x[289], x[281], x[280], x[279], x[278], x[277], x[276], x[230], x[229], x[228], x[227], x[226], x[225], x[29], x[28], x[222], x[221], x[43], x[42], x[41], x[40], x[39], x[38], x[239], x[238], x[26], x[25], x[24], x[23], x[22], x[21], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[205], x[204], x[335], x[291], x[18], x[198], x[195], x[194], x[193], x[192], x[191]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[180], x[163], x[182], x[181], x[95], x[165], x[164], x[265], x[214], x[112], x[282], x[231], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[162], x[161], x[160], x[159], x[158], x[157], x[267], x[266], x[216], x[215], x[44], x[114], x[113], x[284], x[283], x[233], x[232], x[27], x[186], x[185], x[94], x[93], x[92], x[91], x[90], x[89], x[168], x[169], x[264], x[263], x[262], x[261], x[260], x[259], x[213], x[212], x[211], x[210], x[209], x[208], x[46], x[45], x[271], x[270], x[111], x[110], x[109], x[108], x[107], x[106], x[288], x[287], x[281], x[280], x[279], x[278], x[277], x[276], x[230], x[229], x[228], x[227], x[226], x[225], x[29], x[28], x[220], x[219], x[43], x[42], x[41], x[40], x[39], x[38], x[237], x[236], x[26], x[25], x[24], x[23], x[22], x[21], x[203], x[202], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[334], x[291], x[18], x[197], x[195], x[194], x[193], x[192], x[191]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[181], x[164], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[96], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[266], x[215], x[283], x[113], x[232], x[184], x[183], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[166], x[167], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[216], x[214], x[212], x[211], x[210], x[209], x[208], x[45], x[286], x[285], x[284], x[282], x[280], x[279], x[278], x[277], x[276], x[269], x[268], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[28], x[218], x[217], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[235], x[234], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[201], x[200], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[333], x[291], x[18], x[196], x[195], x[194], x[193], x[192], x[191]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[165], x[182], x[164], x[163], x[267], x[181], x[180], x[97], x[216], x[114], x[284], x[233], x[155], x[156], x[162], x[161], x[160], x[159], x[158], x[157], x[266], x[265], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[215], x[214], x[46], x[258], x[257], x[113], x[112], x[275], x[274], x[283], x[282], x[232], x[231], x[29], x[264], x[263], x[262], x[261], x[260], x[259], x[94], x[93], x[92], x[91], x[90], x[89], x[207], x[206], x[213], x[212], x[211], x[210], x[209], x[208], x[45], x[44], x[111], x[110], x[109], x[108], x[107], x[106], x[281], x[280], x[279], x[278], x[277], x[276], x[224], x[223], x[230], x[229], x[228], x[227], x[226], x[225], x[28], x[27], x[43], x[42], x[41], x[40], x[39], x[38], x[26], x[25], x[24], x[23], x[22], x[21], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[190], x[189], x[332], x[291], x[18], x[199], x[195], x[194], x[193], x[192], x[191]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[188], x[187], x[170], x[171], x[205], x[204], x[222], x[221], x[339], x[186], x[185], x[168], x[169], x[203], x[202], x[220], x[219], x[338], x[184], x[183], x[166], x[167], x[201], x[200], x[218], x[217], x[337], x[165], x[182], x[199], x[164], x[163], x[267], x[181], x[180], x[97], x[198], x[197], x[155], x[156], x[162], x[161], x[160], x[159], x[158], x[157], x[266], x[265], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[46], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[264], x[263], x[262], x[261], x[260], x[259], x[94], x[93], x[92], x[91], x[90], x[89], x[45], x[44], x[213], x[43], x[42], x[41], x[40], x[39], x[38], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[207], x[206], x[336], x[291], x[18], x[216], x[212], x[211], x[210], x[209], x[208]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[180], x[163], x[197], x[182], x[181], x[95], x[165], x[164], x[265], x[199], x[198], x[214], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[162], x[161], x[160], x[159], x[158], x[157], x[267], x[266], x[44], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[188], x[187], x[94], x[93], x[92], x[91], x[90], x[89], x[170], x[171], x[264], x[263], x[262], x[261], x[260], x[259], x[46], x[45], x[205], x[204], x[213], x[43], x[42], x[41], x[40], x[39], x[38], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[222], x[221], x[339], x[291], x[18], x[215], x[212], x[211], x[210], x[209], x[208]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[180], x[163], x[197], x[182], x[181], x[95], x[165], x[164], x[265], x[199], x[198], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[162], x[161], x[160], x[159], x[158], x[157], x[267], x[266], x[44], x[196], x[195], x[194], x[193], x[192], x[191], x[216], x[215], x[186], x[185], x[94], x[93], x[92], x[91], x[90], x[89], x[168], x[169], x[264], x[263], x[262], x[261], x[260], x[259], x[46], x[45], x[203], x[202], x[213], x[43], x[42], x[41], x[40], x[39], x[38], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[220], x[219], x[338], x[291], x[18], x[214], x[212], x[211], x[210], x[209], x[208]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[181], x[164], x[198], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[96], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[266], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[215], x[184], x[183], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[166], x[167], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[45], x[201], x[200], x[216], x[214], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[218], x[217], x[337], x[291], x[18], x[213], x[212], x[211], x[210], x[209], x[208]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[165], x[182], x[199], x[164], x[163], x[267], x[181], x[180], x[97], x[198], x[197], x[155], x[156], x[162], x[161], x[160], x[159], x[158], x[157], x[266], x[265], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[46], x[190], x[189], x[196], x[195], x[194], x[193], x[192], x[191], x[215], x[214], x[264], x[263], x[262], x[261], x[260], x[259], x[94], x[93], x[92], x[91], x[90], x[89], x[45], x[44], x[213], x[43], x[42], x[41], x[40], x[39], x[38], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[207], x[206], x[336], x[291], x[18], x[216], x[212], x[211], x[210], x[209], x[208]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[273], x[272], x[290], x[289], x[119], x[120], x[102], x[103], x[256], x[255], x[153], x[154], x[239], x[238], x[343], x[232], x[271], x[270], x[288], x[287], x[117], x[118], x[100], x[101], x[254], x[253], x[151], x[152], x[237], x[236], x[342], x[231], x[286], x[285], x[269], x[268], x[115], x[116], x[98], x[99], x[252], x[251], x[149], x[150], x[235], x[234], x[341], x[230], x[267], x[97], x[266], x[265], x[114], x[284], x[250], x[96], x[95], x[182], x[80], x[148], x[258], x[257], x[264], x[263], x[262], x[261], x[260], x[259], x[113], x[112], x[275], x[274], x[283], x[282], x[249], x[248], x[199], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[104], x[105], x[79], x[78], x[147], x[146], x[131], x[111], x[110], x[109], x[108], x[107], x[106], x[281], x[280], x[279], x[278], x[277], x[276], x[241], x[240], x[247], x[246], x[245], x[244], x[243], x[242], x[198], x[197], x[179], x[178], x[177], x[176], x[175], x[174], x[77], x[76], x[75], x[74], x[73], x[72], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[196], x[195], x[194], x[193], x[192], x[191], x[128], x[127], x[126], x[125], x[124], x[123], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[224], x[223], x[340], x[291], x[18], x[233], x[229], x[228], x[227], x[226], x[225]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[265], x[95], x[267], x[266], x[112], x[282], x[248], x[78], x[97], x[96], x[180], x[146], x[264], x[263], x[262], x[261], x[260], x[259], x[114], x[113], x[284], x[283], x[250], x[249], x[197], x[80], x[79], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[148], x[147], x[129], x[273], x[272], x[111], x[110], x[109], x[108], x[107], x[106], x[290], x[289], x[281], x[280], x[279], x[278], x[277], x[276], x[247], x[246], x[245], x[244], x[243], x[242], x[199], x[198], x[119], x[120], x[77], x[76], x[75], x[74], x[73], x[72], x[102], x[103], x[179], x[178], x[177], x[176], x[175], x[174], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[256], x[255], x[196], x[195], x[194], x[193], x[192], x[191], x[153], x[154], x[128], x[127], x[126], x[125], x[124], x[123], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[239], x[238], x[343], x[291], x[18], x[232], x[229], x[228], x[227], x[226], x[225]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[265], x[95], x[267], x[266], x[112], x[282], x[248], x[78], x[97], x[96], x[180], x[146], x[264], x[263], x[262], x[261], x[260], x[259], x[114], x[113], x[284], x[283], x[250], x[249], x[197], x[80], x[79], x[94], x[93], x[92], x[91], x[90], x[89], x[182], x[181], x[148], x[147], x[129], x[271], x[270], x[111], x[110], x[109], x[108], x[107], x[106], x[288], x[287], x[281], x[280], x[279], x[278], x[277], x[276], x[247], x[246], x[245], x[244], x[243], x[242], x[199], x[198], x[117], x[118], x[77], x[76], x[75], x[74], x[73], x[72], x[100], x[101], x[179], x[178], x[177], x[176], x[175], x[174], x[145], x[144], x[143], x[142], x[141], x[140], x[131], x[130], x[254], x[253], x[196], x[195], x[194], x[193], x[192], x[191], x[151], x[152], x[128], x[127], x[126], x[125], x[124], x[123], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[237], x[236], x[342], x[291], x[18], x[231], x[229], x[228], x[227], x[226], x[225]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[266], x[96], x[283], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[113], x[249], x[79], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[181], x[147], x[286], x[285], x[284], x[282], x[280], x[279], x[278], x[277], x[276], x[269], x[268], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[198], x[115], x[116], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[98], x[99], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[130], x[252], x[251], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[149], x[150], x[131], x[129], x[127], x[126], x[125], x[124], x[123], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[235], x[234], x[341], x[291], x[18], x[230], x[229], x[228], x[227], x[226], x[225]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[267], x[97], x[266], x[265], x[114], x[284], x[250], x[96], x[95], x[182], x[80], x[148], x[258], x[257], x[264], x[263], x[262], x[261], x[260], x[259], x[113], x[112], x[275], x[274], x[283], x[282], x[249], x[248], x[199], x[87], x[88], x[94], x[93], x[92], x[91], x[90], x[89], x[181], x[180], x[104], x[105], x[79], x[78], x[147], x[146], x[131], x[111], x[110], x[109], x[108], x[107], x[106], x[281], x[280], x[279], x[278], x[277], x[276], x[241], x[240], x[247], x[246], x[245], x[244], x[243], x[242], x[198], x[197], x[179], x[178], x[177], x[176], x[175], x[174], x[77], x[76], x[75], x[74], x[73], x[72], x[138], x[139], x[145], x[144], x[143], x[142], x[141], x[140], x[130], x[129], x[196], x[195], x[194], x[193], x[192], x[191], x[128], x[127], x[126], x[125], x[124], x[123], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[224], x[223], x[340], x[291], x[18], x[233], x[229], x[228], x[227], x[226], x[225]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[273], x[272], x[290], x[289], x[68], x[69], x[85], x[86], x[239], x[238], x[34], x[35], x[256], x[255], x[347], x[249], x[271], x[270], x[288], x[287], x[66], x[67], x[83], x[84], x[237], x[236], x[32], x[33], x[254], x[253], x[346], x[248], x[286], x[285], x[269], x[268], x[81], x[82], x[65], x[64], x[235], x[234], x[30], x[31], x[252], x[251], x[345], x[247], x[267], x[80], x[266], x[265], x[114], x[284], x[233], x[63], x[79], x[78], x[165], x[258], x[257], x[264], x[263], x[262], x[261], x[260], x[259], x[113], x[112], x[275], x[274], x[283], x[282], x[232], x[231], x[29], x[54], x[53], x[62], x[61], x[70], x[71], x[77], x[76], x[75], x[74], x[73], x[72], x[164], x[163], x[148], x[111], x[110], x[109], x[108], x[107], x[106], x[281], x[280], x[279], x[278], x[277], x[276], x[224], x[223], x[230], x[229], x[228], x[227], x[226], x[225], x[28], x[27], x[60], x[59], x[58], x[57], x[56], x[55], x[162], x[161], x[160], x[159], x[158], x[157], x[19], x[20], x[147], x[146], x[26], x[25], x[24], x[23], x[22], x[21], x[145], x[144], x[143], x[142], x[141], x[140], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[241], x[240], x[344], x[291], x[18], x[250], x[246], x[245], x[244], x[243], x[242]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[265], x[78], x[267], x[266], x[112], x[282], x[231], x[61], x[80], x[79], x[163], x[264], x[263], x[262], x[261], x[260], x[259], x[114], x[113], x[284], x[283], x[233], x[232], x[27], x[63], x[62], x[77], x[76], x[75], x[74], x[73], x[72], x[165], x[164], x[146], x[273], x[272], x[111], x[110], x[109], x[108], x[107], x[106], x[290], x[289], x[281], x[280], x[279], x[278], x[277], x[276], x[230], x[229], x[228], x[227], x[226], x[225], x[29], x[28], x[68], x[69], x[60], x[59], x[58], x[57], x[56], x[55], x[85], x[86], x[162], x[161], x[160], x[159], x[158], x[157], x[148], x[147], x[239], x[238], x[26], x[25], x[24], x[23], x[22], x[21], x[34], x[35], x[145], x[144], x[143], x[142], x[141], x[140], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[256], x[255], x[347], x[291], x[18], x[249], x[246], x[245], x[244], x[243], x[242]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[265], x[78], x[267], x[266], x[112], x[282], x[231], x[61], x[80], x[79], x[163], x[264], x[263], x[262], x[261], x[260], x[259], x[114], x[113], x[284], x[283], x[233], x[232], x[27], x[63], x[62], x[77], x[76], x[75], x[74], x[73], x[72], x[165], x[164], x[146], x[271], x[270], x[111], x[110], x[109], x[108], x[107], x[106], x[288], x[287], x[281], x[280], x[279], x[278], x[277], x[276], x[230], x[229], x[228], x[227], x[226], x[225], x[29], x[28], x[66], x[67], x[60], x[59], x[58], x[57], x[56], x[55], x[83], x[84], x[162], x[161], x[160], x[159], x[158], x[157], x[148], x[147], x[237], x[236], x[26], x[25], x[24], x[23], x[22], x[21], x[32], x[33], x[145], x[144], x[143], x[142], x[141], x[140], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[254], x[253], x[346], x[291], x[18], x[248], x[246], x[245], x[244], x[243], x[242]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[266], x[79], x[283], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[113], x[232], x[80], x[78], x[76], x[75], x[74], x[73], x[72], x[164], x[62], x[286], x[285], x[284], x[282], x[280], x[279], x[278], x[277], x[276], x[269], x[268], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[28], x[81], x[82], x[165], x[163], x[161], x[160], x[159], x[158], x[157], x[65], x[64], x[63], x[61], x[59], x[58], x[57], x[56], x[55], x[147], x[235], x[234], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[30], x[31], x[148], x[146], x[144], x[143], x[142], x[141], x[140], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[252], x[251], x[345], x[291], x[18], x[247], x[246], x[245], x[244], x[243], x[242]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[267], x[80], x[266], x[265], x[114], x[284], x[233], x[63], x[79], x[78], x[165], x[258], x[257], x[264], x[263], x[262], x[261], x[260], x[259], x[113], x[112], x[275], x[274], x[283], x[282], x[232], x[231], x[29], x[54], x[53], x[62], x[61], x[70], x[71], x[77], x[76], x[75], x[74], x[73], x[72], x[164], x[163], x[148], x[111], x[110], x[109], x[108], x[107], x[106], x[281], x[280], x[279], x[278], x[277], x[276], x[224], x[223], x[230], x[229], x[228], x[227], x[226], x[225], x[28], x[27], x[60], x[59], x[58], x[57], x[56], x[55], x[162], x[161], x[160], x[159], x[158], x[157], x[19], x[20], x[147], x[146], x[26], x[25], x[24], x[23], x[22], x[21], x[145], x[144], x[143], x[142], x[141], x[140], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[241], x[240], x[344], x[291], x[18], x[250], x[246], x[245], x[244], x[243], x[242]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[256], x[255], x[239], x[238], x[205], x[204], x[222], x[221], x[290], x[289], x[188], x[187], x[273], x[272], x[351], x[266], x[254], x[253], x[237], x[236], x[203], x[202], x[220], x[219], x[288], x[287], x[186], x[185], x[271], x[270], x[350], x[265], x[252], x[251], x[235], x[234], x[218], x[217], x[201], x[200], x[286], x[285], x[184], x[183], x[269], x[268], x[349], x[264], x[233], x[250], x[232], x[231], x[29], x[249], x[248], x[199], x[216], x[46], x[182], x[224], x[223], x[230], x[229], x[228], x[227], x[226], x[225], x[28], x[27], x[241], x[240], x[247], x[246], x[245], x[244], x[243], x[242], x[198], x[197], x[284], x[190], x[189], x[215], x[214], x[207], x[206], x[45], x[44], x[181], x[180], x[97], x[26], x[25], x[24], x[23], x[22], x[21], x[196], x[195], x[194], x[193], x[192], x[191], x[275], x[274], x[283], x[282], x[213], x[212], x[211], x[210], x[209], x[208], x[43], x[42], x[41], x[40], x[39], x[38], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[281], x[280], x[279], x[278], x[277], x[276], x[94], x[93], x[92], x[91], x[90], x[89], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[258], x[257], x[348], x[291], x[18], x[267], x[263], x[262], x[261], x[260], x[259]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[248], x[231], x[250], x[249], x[197], x[233], x[232], x[27], x[214], x[44], x[180], x[247], x[246], x[245], x[244], x[243], x[242], x[199], x[198], x[230], x[229], x[228], x[227], x[226], x[225], x[29], x[28], x[282], x[216], x[215], x[46], x[45], x[182], x[181], x[95], x[256], x[255], x[196], x[195], x[194], x[193], x[192], x[191], x[239], x[238], x[26], x[25], x[24], x[23], x[22], x[21], x[284], x[283], x[205], x[204], x[213], x[212], x[211], x[210], x[209], x[208], x[222], x[221], x[43], x[42], x[41], x[40], x[39], x[38], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[290], x[289], x[281], x[280], x[279], x[278], x[277], x[276], x[188], x[187], x[94], x[93], x[92], x[91], x[90], x[89], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[273], x[272], x[351], x[291], x[18], x[266], x[263], x[262], x[261], x[260], x[259]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[248], x[231], x[250], x[249], x[197], x[233], x[232], x[27], x[214], x[44], x[180], x[247], x[246], x[245], x[244], x[243], x[242], x[199], x[198], x[230], x[229], x[228], x[227], x[226], x[225], x[29], x[28], x[282], x[216], x[215], x[46], x[45], x[182], x[181], x[95], x[254], x[253], x[196], x[195], x[194], x[193], x[192], x[191], x[237], x[236], x[26], x[25], x[24], x[23], x[22], x[21], x[284], x[283], x[203], x[202], x[213], x[212], x[211], x[210], x[209], x[208], x[220], x[219], x[43], x[42], x[41], x[40], x[39], x[38], x[179], x[178], x[177], x[176], x[175], x[174], x[97], x[96], x[288], x[287], x[281], x[280], x[279], x[278], x[277], x[276], x[186], x[185], x[94], x[93], x[92], x[91], x[90], x[89], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[271], x[270], x[350], x[291], x[18], x[265], x[263], x[262], x[261], x[260], x[259]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[249], x[232], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[198], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[28], x[45], x[215], x[181], x[252], x[251], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[235], x[234], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[283], x[218], x[217], x[46], x[44], x[42], x[41], x[40], x[39], x[38], x[201], x[200], x[216], x[214], x[212], x[211], x[210], x[209], x[208], x[182], x[180], x[178], x[177], x[176], x[175], x[174], x[96], x[286], x[285], x[284], x[282], x[280], x[279], x[278], x[277], x[276], x[184], x[183], x[97], x[95], x[93], x[92], x[91], x[90], x[89], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[269], x[268], x[349], x[291], x[18], x[264], x[263], x[262], x[261], x[260], x[259]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[233], x[250], x[232], x[231], x[29], x[249], x[248], x[199], x[216], x[46], x[182], x[224], x[223], x[230], x[229], x[228], x[227], x[226], x[225], x[28], x[27], x[241], x[240], x[247], x[246], x[245], x[244], x[243], x[242], x[198], x[197], x[284], x[190], x[189], x[215], x[214], x[207], x[206], x[45], x[44], x[181], x[180], x[97], x[26], x[25], x[24], x[23], x[22], x[21], x[196], x[195], x[194], x[193], x[192], x[191], x[275], x[274], x[283], x[282], x[213], x[212], x[211], x[210], x[209], x[208], x[43], x[42], x[41], x[40], x[39], x[38], x[173], x[172], x[179], x[178], x[177], x[176], x[175], x[174], x[96], x[95], x[281], x[280], x[279], x[278], x[277], x[276], x[94], x[93], x[92], x[91], x[90], x[89], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[258], x[257], x[348], x[291], x[18], x[267], x[263], x[262], x[261], x[260], x[259]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[256], x[255], x[239], x[238], x[273], x[272], x[290], x[289], x[355], x[283], x[254], x[253], x[237], x[236], x[271], x[270], x[288], x[287], x[354], x[282], x[252], x[251], x[235], x[234], x[269], x[268], x[286], x[285], x[353], x[281], x[233], x[250], x[232], x[231], x[29], x[249], x[248], x[199], x[267], x[224], x[223], x[230], x[229], x[228], x[227], x[226], x[225], x[28], x[27], x[241], x[240], x[247], x[246], x[245], x[244], x[243], x[242], x[198], x[197], x[266], x[265], x[114], x[26], x[25], x[24], x[23], x[22], x[21], x[196], x[195], x[194], x[193], x[192], x[191], x[258], x[257], x[264], x[263], x[262], x[261], x[260], x[259], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[275], x[274], x[352], x[291], x[18], x[284], x[280], x[279], x[278], x[277], x[276]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[248], x[231], x[250], x[249], x[197], x[233], x[232], x[27], x[265], x[247], x[246], x[245], x[244], x[243], x[242], x[199], x[198], x[230], x[229], x[228], x[227], x[226], x[225], x[29], x[28], x[267], x[266], x[112], x[256], x[255], x[196], x[195], x[194], x[193], x[192], x[191], x[239], x[238], x[26], x[25], x[24], x[23], x[22], x[21], x[264], x[263], x[262], x[261], x[260], x[259], x[114], x[113], x[273], x[272], x[111], x[110], x[109], x[108], x[107], x[106], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[290], x[289], x[355], x[291], x[18], x[283], x[280], x[279], x[278], x[277], x[276]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[248], x[231], x[250], x[249], x[197], x[233], x[232], x[27], x[265], x[247], x[246], x[245], x[244], x[243], x[242], x[199], x[198], x[230], x[229], x[228], x[227], x[226], x[225], x[29], x[28], x[267], x[266], x[112], x[254], x[253], x[196], x[195], x[194], x[193], x[192], x[191], x[237], x[236], x[26], x[25], x[24], x[23], x[22], x[21], x[264], x[263], x[262], x[261], x[260], x[259], x[114], x[113], x[271], x[270], x[111], x[110], x[109], x[108], x[107], x[106], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[288], x[287], x[354], x[291], x[18], x[282], x[280], x[279], x[278], x[277], x[276]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[249], x[232], x[250], x[248], x[246], x[245], x[244], x[243], x[242], x[198], x[233], x[231], x[229], x[228], x[227], x[226], x[225], x[28], x[266], x[252], x[251], x[199], x[197], x[195], x[194], x[193], x[192], x[191], x[235], x[234], x[29], x[27], x[25], x[24], x[23], x[22], x[21], x[267], x[265], x[263], x[262], x[261], x[260], x[259], x[113], x[269], x[268], x[114], x[112], x[110], x[109], x[108], x[107], x[106], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[286], x[285], x[353], x[291], x[18], x[281], x[280], x[279], x[278], x[277], x[276]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[233], x[250], x[232], x[231], x[29], x[249], x[248], x[199], x[267], x[224], x[223], x[230], x[229], x[228], x[227], x[226], x[225], x[28], x[27], x[241], x[240], x[247], x[246], x[245], x[244], x[243], x[242], x[198], x[197], x[266], x[265], x[114], x[26], x[25], x[24], x[23], x[22], x[21], x[196], x[195], x[194], x[193], x[192], x[191], x[258], x[257], x[264], x[263], x[262], x[261], x[260], x[259], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[275], x[274], x[352], x[291], x[18], x[284], x[280], x[279], x[278], x[277], x[276]}), .y(y[189]));
endmodule

